-- This file was generated with hex2rom written by Daniel Wallner

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ProgramROM is
    port(
        A   : in std_logic_vector(13 downto 0);
        D   : out std_logic_vector(7 downto 0)
    );
end ProgramROM;

architecture rtl of ProgramROM is
    subtype ROM_WORD is std_logic_vector(7 downto 0);
    type ROM_TABLE is array(0 to 16383) of ROM_WORD;
    constant ROM: ROM_TABLE := ROM_TABLE'(
        "00000010", -- 0x0000
        "00000000", -- 0x0001
        "00011110", -- 0x0002
        "00000010", -- 0x0003
        "00010110", -- 0x0004
        "01111100", -- 0x0005
        "00010010", -- 0x0006
        "00100100", -- 0x0007
        "10010101", -- 0x0008
        "00010010", -- 0x0009
        "00100001", -- 0x000A
        "10100100", -- 0x000B
        "00010010", -- 0x000C
        "00011001", -- 0x000D
        "01001000", -- 0x000E
        "00010010", -- 0x000F
        "00011111", -- 0x0010
        "00001000", -- 0x0011
        "00100010", -- 0x0012
        "00000010", -- 0x0013
        "00011110", -- 0x0014
        "00010011", -- 0x0015
        "00010010", -- 0x0016
        "00100100", -- 0x0017
        "01110011", -- 0x0018
        "01001000", -- 0x0019
        "00100010", -- 0x001A
        "00000010", -- 0x001B
        "00010001", -- 0x001C
        "10000000", -- 0x001D
        "01110101", -- 0x001E
        "11010000", -- 0x001F
        "00000000", -- 0x0020
        "01110101", -- 0x0021
        "10011111", -- 0x0022
        "00000000", -- 0x0023
        "01110101", -- 0x0024
        "10001111", -- 0x0025
        "10000000", -- 0x0026
        "01110101", -- 0x0027
        "10000001", -- 0x0028
        "00100000", -- 0x0029
        "00010010", -- 0x002A
        "00000110", -- 0x002B
        "01100000", -- 0x002C
        "11100100", -- 0x002D
        "11111111", -- 0x002E
        "11111110", -- 0x002F
        "00010010", -- 0x0030
        "00001011", -- 0x0031
        "11101111", -- 0x0032
        "00010010", -- 0x0033
        "00100100", -- 0x0034
        "10100000", -- 0x0035
        "00110010", -- 0x0036
        "00000000", -- 0x0037
        "00000001", -- 0x0038
        "00000000", -- 0x0039
        "00000000", -- 0x003A
        "00000000", -- 0x003B
        "00000000", -- 0x003C
        "00100111", -- 0x003D
        "00010000", -- 0x003E
        "00000000", -- 0x003F
        "00000000", -- 0x0040
        "00000000", -- 0x0041
        "00000000", -- 0x0042
        "00000000", -- 0x0043
        "00000000", -- 0x0044
        "00000000", -- 0x0045
        "00000000", -- 0x0046
        "00000000", -- 0x0047
        "11111111", -- 0x0048
        "00000000", -- 0x0049
        "00000000", -- 0x004A
        "00000000", -- 0x004B
        "00000000", -- 0x004C
        "00000000", -- 0x004D
        "00000000", -- 0x004E
        "10100000", -- 0x004F
        "10100000", -- 0x0050
        "10100000", -- 0x0051
        "10100000", -- 0x0052
        "10100000", -- 0x0053
        "10100000", -- 0x0054
        "10100000", -- 0x0055
        "10100000", -- 0x0056
        "10100000", -- 0x0057
        "10100000", -- 0x0058
        "10100000", -- 0x0059
        "10100000", -- 0x005A
        "10100000", -- 0x005B
        "10100000", -- 0x005C
        "10100000", -- 0x005D
        "10100000", -- 0x005E
        "10100000", -- 0x005F
        "10100000", -- 0x0060
        "10100000", -- 0x0061
        "10100000", -- 0x0062
        "10011111", -- 0x0063
        "10011111", -- 0x0064
        "10011110", -- 0x0065
        "10011110", -- 0x0066
        "10011101", -- 0x0067
        "10011101", -- 0x0068
        "10011100", -- 0x0069
        "10011100", -- 0x006A
        "10011011", -- 0x006B
        "10011010", -- 0x006C
        "10011010", -- 0x006D
        "10011001", -- 0x006E
        "10011001", -- 0x006F
        "10011000", -- 0x0070
        "10011000", -- 0x0071
        "10010111", -- 0x0072
        "10010111", -- 0x0073
        "10010110", -- 0x0074
        "10010101", -- 0x0075
        "10010011", -- 0x0076
        "10010010", -- 0x0077
        "10010001", -- 0x0078
        "10010000", -- 0x0079
        "10010000", -- 0x007A
        "10001111", -- 0x007B
        "10001110", -- 0x007C
        "10001110", -- 0x007D
        "10001101", -- 0x007E
        "10001101", -- 0x007F
        "10001100", -- 0x0080
        "10001011", -- 0x0081
        "10001010", -- 0x0082
        "10001001", -- 0x0083
        "10001000", -- 0x0084
        "10000111", -- 0x0085
        "10000110", -- 0x0086
        "10000110", -- 0x0087
        "10000101", -- 0x0088
        "10000101", -- 0x0089
        "10000100", -- 0x008A
        "10000100", -- 0x008B
        "10000011", -- 0x008C
        "10000011", -- 0x008D
        "10000010", -- 0x008E
        "10000001", -- 0x008F
        "10000000", -- 0x0090
        "01111111", -- 0x0091
        "01111111", -- 0x0092
        "01111110", -- 0x0093
        "01111101", -- 0x0094
        "01111100", -- 0x0095
        "01111011", -- 0x0096
        "01111010", -- 0x0097
        "01111001", -- 0x0098
        "01111000", -- 0x0099
        "01110111", -- 0x009A
        "01110111", -- 0x009B
        "01110110", -- 0x009C
        "01110101", -- 0x009D
        "01110101", -- 0x009E
        "01110100", -- 0x009F
        "01110100", -- 0x00A0
        "01101110", -- 0x00A1
        "01101110", -- 0x00A2
        "01101101", -- 0x00A3
        "01101101", -- 0x00A4
        "01101101", -- 0x00A5
        "01101101", -- 0x00A6
        "01101100", -- 0x00A7
        "01101100", -- 0x00A8
        "01101100", -- 0x00A9
        "01101011", -- 0x00AA
        "01101011", -- 0x00AB
        "01101011", -- 0x00AC
        "01101010", -- 0x00AD
        "01101010", -- 0x00AE
        "01101010", -- 0x00AF
        "01101010", -- 0x00B0
        "01101001", -- 0x00B1
        "01101001", -- 0x00B2
        "01100111", -- 0x00B3
        "01100110", -- 0x00B4
        "01100100", -- 0x00B5
        "01100011", -- 0x00B6
        "01100011", -- 0x00B7
        "01100010", -- 0x00B8
        "01100010", -- 0x00B9
        "01100001", -- 0x00BA
        "01100001", -- 0x00BB
        "01100000", -- 0x00BC
        "01100000", -- 0x00BD
        "01011111", -- 0x00BE
        "01011110", -- 0x00BF
        "01011110", -- 0x00C0
        "01011101", -- 0x00C1
        "01011101", -- 0x00C2
        "01011100", -- 0x00C3
        "01011100", -- 0x00C4
        "01011011", -- 0x00C5
        "01011011", -- 0x00C6
        "01011010", -- 0x00C7
        "01011001", -- 0x00C8
        "01011001", -- 0x00C9
        "01011000", -- 0x00CA
        "01011000", -- 0x00CB
        "01010111", -- 0x00CC
        "01010111", -- 0x00CD
        "01010110", -- 0x00CE
        "01010110", -- 0x00CF
        "01010101", -- 0x00D0
        "01010101", -- 0x00D1
        "01010100", -- 0x00D2
        "01010011", -- 0x00D3
        "01010010", -- 0x00D4
        "01010001", -- 0x00D5
        "01010000", -- 0x00D6
        "01001111", -- 0x00D7
        "01001111", -- 0x00D8
        "01001110", -- 0x00D9
        "01001110", -- 0x00DA
        "01001101", -- 0x00DB
        "01001101", -- 0x00DC
        "01001100", -- 0x00DD
        "01001100", -- 0x00DE
        "01001011", -- 0x00DF
        "01001010", -- 0x00E0
        "01001001", -- 0x00E1
        "01001000", -- 0x00E2
        "01001000", -- 0x00E3
        "01000111", -- 0x00E4
        "01000110", -- 0x00E5
        "01000101", -- 0x00E6
        "01000101", -- 0x00E7
        "01000100", -- 0x00E8
        "01000011", -- 0x00E9
        "01000010", -- 0x00EA
        "01000010", -- 0x00EB
        "01000001", -- 0x00EC
        "01000000", -- 0x00ED
        "00111111", -- 0x00EE
        "00111110", -- 0x00EF
        "00111110", -- 0x00F0
        "00111101", -- 0x00F1
        "00111100", -- 0x00F2
        "00111011", -- 0x00F3
        "00111010", -- 0x00F4
        "00111001", -- 0x00F5
        "00111000", -- 0x00F6
        "00110111", -- 0x00F7
        "00110110", -- 0x00F8
        "00110101", -- 0x00F9
        "00110100", -- 0x00FA
        "00110100", -- 0x00FB
        "00110011", -- 0x00FC
        "00110010", -- 0x00FD
        "00110001", -- 0x00FE
        "00110000", -- 0x00FF
        "00101111", -- 0x0100
        "00101111", -- 0x0101
        "00101110", -- 0x0102
        "00101101", -- 0x0103
        "00101100", -- 0x0104
        "00101011", -- 0x0105
        "00101010", -- 0x0106
        "00101001", -- 0x0107
        "00101000", -- 0x0108
        "00100111", -- 0x0109
        "00100110", -- 0x010A
        "00100101", -- 0x010B
        "00100101", -- 0x010C
        "00100100", -- 0x010D
        "00100011", -- 0x010E
        "00100010", -- 0x010F
        "00100010", -- 0x0110
        "00100001", -- 0x0111
        "00100001", -- 0x0112
        "00100000", -- 0x0113
        "00100000", -- 0x0114
        "00011111", -- 0x0115
        "00011111", -- 0x0116
        "00011110", -- 0x0117
        "00011101", -- 0x0118
        "00011100", -- 0x0119
        "00011011", -- 0x011A
        "00011010", -- 0x011B
        "00011001", -- 0x011C
        "00011001", -- 0x011D
        "00011000", -- 0x011E
        "00011000", -- 0x011F
        "00010111", -- 0x0120
        "00010111", -- 0x0121
        "00010110", -- 0x0122
        "00010110", -- 0x0123
        "00010110", -- 0x0124
        "00010101", -- 0x0125
        "00010101", -- 0x0126
        "00010100", -- 0x0127
        "00010100", -- 0x0128
        "00010011", -- 0x0129
        "00010010", -- 0x012A
        "00010001", -- 0x012B
        "00010001", -- 0x012C
        "00010000", -- 0x012D
        "00001111", -- 0x012E
        "00001101", -- 0x012F
        "00001100", -- 0x0130
        "00001010", -- 0x0131
        "00001001", -- 0x0132
        "00001000", -- 0x0133
        "00000111", -- 0x0134
        "00000111", -- 0x0135
        "00000110", -- 0x0136
        "00000101", -- 0x0137
        "00000100", -- 0x0138
        "00000011", -- 0x0139
        "00000010", -- 0x013A
        "00000001", -- 0x013B
        "00000000", -- 0x013C
        "00000000", -- 0x013D
        "00000000", -- 0x013E
        "00000000", -- 0x013F
        "00000000", -- 0x0140
        "00000000", -- 0x0141
        "00000000", -- 0x0142
        "00000000", -- 0x0143
        "00000000", -- 0x0144
        "00000000", -- 0x0145
        "00000000", -- 0x0146
        "00000000", -- 0x0147
        "00000000", -- 0x0148
        "00000000", -- 0x0149
        "00000000", -- 0x014A
        "00000000", -- 0x014B
        "00000000", -- 0x014C
        "00000000", -- 0x014D
        "00000000", -- 0x014E
        "10001111", -- 0x014F
        "00001100", -- 0x0150
        "10001110", -- 0x0151
        "00001011", -- 0x0152
        "00010010", -- 0x0153
        "00011001", -- 0x0154
        "01001000", -- 0x0155
        "10010000", -- 0x0156
        "00000001", -- 0x0157
        "10011001", -- 0x0158
        "00010010", -- 0x0159
        "00100001", -- 0x015A
        "11001000", -- 0x015B
        "10000101", -- 0x015C
        "00001100", -- 0x015D
        "00001110", -- 0x015E
        "10000101", -- 0x015F
        "00001011", -- 0x0160
        "00001101", -- 0x0161
        "00000101", -- 0x0162
        "00001110", -- 0x0163
        "11100101", -- 0x0164
        "00001110", -- 0x0165
        "01110000", -- 0x0166
        "00000010", -- 0x0167
        "00000101", -- 0x0168
        "00001101", -- 0x0169
        "10101101", -- 0x016A
        "00001110", -- 0x016B
        "10101100", -- 0x016C
        "00001101", -- 0x016D
        "01111010", -- 0x016E
        "00000000", -- 0x016F
        "01111011", -- 0x0170
        "00000011", -- 0x0171
        "01111110", -- 0x0172
        "00000001", -- 0x0173
        "01111111", -- 0x0174
        "10011110", -- 0x0175
        "00010010", -- 0x0176
        "00010100", -- 0x0177
        "01111001", -- 0x0178
        "10010000", -- 0x0179
        "00000001", -- 0x017A
        "10011101", -- 0x017B
        "11100000", -- 0x017C
        "00000100", -- 0x017D
        "11110000", -- 0x017E
        "01111000", -- 0x017F
        "11001100", -- 0x0180
        "10000101", -- 0x0181
        "00001110", -- 0x0182
        "10000010", -- 0x0183
        "10000101", -- 0x0184
        "00001101", -- 0x0185
        "10000011", -- 0x0186
        "11100000", -- 0x0187
        "10010000", -- 0x0188
        "00011001", -- 0x0189
        "10111010", -- 0x018A
        "01110101", -- 0x018B
        "11110000", -- 0x018C
        "00010011", -- 0x018D
        "00010010", -- 0x018E
        "00011011", -- 0x018F
        "11110111", -- 0x0190
        "00000010", -- 0x0191
        "00000011", -- 0x0192
        "00101000", -- 0x0193
        "11100101", -- 0x0194
        "00001100", -- 0x0195
        "00100100", -- 0x0196
        "00000010", -- 0x0197
        "11111001", -- 0x0198
        "11100100", -- 0x0199
        "00110101", -- 0x019A
        "00001011", -- 0x019B
        "00010010", -- 0x019C
        "00100100", -- 0x019D
        "10011001", -- 0x019E
        "10010000", -- 0x019F
        "00010111", -- 0x01A0
        "11010000", -- 0x01A1
        "00010010", -- 0x01A2
        "00100001", -- 0x01A3
        "01101000", -- 0x01A4
        "10010000", -- 0x01A5
        "00010111", -- 0x01A6
        "11010001", -- 0x01A7
        "11110000", -- 0x01A8
        "01111100", -- 0x01A9
        "00000000", -- 0x01AA
        "01111101", -- 0x01AB
        "00000010", -- 0x01AC
        "01111110", -- 0x01AD
        "00010111", -- 0x01AE
        "01111111", -- 0x01AF
        "11010000", -- 0x01B0
        "00010010", -- 0x01B1
        "00010111", -- 0x01B2
        "10001110", -- 0x01B3
        "10010000", -- 0x01B4
        "00010111", -- 0x01B5
        "11010010", -- 0x01B6
        "11110000", -- 0x01B7
        "01111110", -- 0x01B8
        "00010111", -- 0x01B9
        "01111111", -- 0x01BA
        "11010000", -- 0x01BB
        "00010010", -- 0x01BC
        "00001101", -- 0x01BD
        "01010011", -- 0x01BE
        "01111000", -- 0x01BF
        "11111111", -- 0x01C0
        "00000010", -- 0x01C1
        "00000011", -- 0x01C2
        "00101000", -- 0x01C3
        "00010010", -- 0x01C4
        "00100000", -- 0x01C5
        "01101000", -- 0x01C6
        "10010000", -- 0x01C7
        "00000001", -- 0x01C8
        "00111110", -- 0x01C9
        "00010010", -- 0x01CA
        "00100100", -- 0x01CB
        "01010100", -- 0x01CC
        "10010000", -- 0x01CD
        "00000001", -- 0x01CE
        "00111110", -- 0x01CF
        "00010010", -- 0x01D0
        "00011111", -- 0x01D1
        "01000100", -- 0x01D2
        "10010000", -- 0x01D3
        "00000001", -- 0x01D4
        "00111110", -- 0x01D5
        "00010010", -- 0x01D6
        "00011111", -- 0x01D7
        "10010001", -- 0x01D8
        "01111000", -- 0x01D9
        "00000000", -- 0x01DA
        "00000010", -- 0x01DB
        "00000011", -- 0x01DC
        "00101000", -- 0x01DD
        "00010010", -- 0x01DE
        "00011111", -- 0x01DF
        "11111001", -- 0x01E0
        "01110100", -- 0x01E1
        "10100000", -- 0x01E2
        "11000011", -- 0x01E3
        "10011001", -- 0x01E4
        "01010000", -- 0x01E5
        "00000011", -- 0x01E6
        "00000010", -- 0x01E7
        "00000011", -- 0x01E8
        "00101000", -- 0x01E9
        "10010000", -- 0x01EA
        "00000001", -- 0x01EB
        "00111101", -- 0x01EC
        "11101001", -- 0x01ED
        "11110000", -- 0x01EE
        "10000000", -- 0x01EF
        "11101000", -- 0x01F0
        "00010010", -- 0x01F1
        "00100001", -- 0x01F2
        "11110110", -- 0x01F3
        "10010000", -- 0x01F4
        "00000001", -- 0x01F5
        "01000011", -- 0x01F6
        "11110000", -- 0x01F7
        "10000000", -- 0x01F8
        "11011111", -- 0x01F9
        "10010000", -- 0x01FA
        "00000001", -- 0x01FB
        "10010110", -- 0x01FC
        "11100000", -- 0x01FD
        "10010000", -- 0x01FE
        "00000001", -- 0x01FF
        "01000101", -- 0x0200
        "11110000", -- 0x0201
        "10000000", -- 0x0202
        "11010101", -- 0x0203
        "00010010", -- 0x0204
        "00100000", -- 0x0205
        "01101000", -- 0x0206
        "10010000", -- 0x0207
        "00000001", -- 0x0208
        "01000000", -- 0x0209
        "00010010", -- 0x020A
        "00100100", -- 0x020B
        "01010100", -- 0x020C
        "10010000", -- 0x020D
        "00000001", -- 0x020E
        "01000000", -- 0x020F
        "00010010", -- 0x0210
        "00011111", -- 0x0211
        "01000100", -- 0x0212
        "10010000", -- 0x0213
        "00000001", -- 0x0214
        "01000000", -- 0x0215
        "10000000", -- 0x0216
        "10111110", -- 0x0217
        "00010010", -- 0x0218
        "00011111", -- 0x0219
        "11111001", -- 0x021A
        "01100100", -- 0x021B
        "00000001", -- 0x021C
        "01100000", -- 0x021D
        "00000110", -- 0x021E
        "11101001", -- 0x021F
        "01100000", -- 0x0220
        "00000011", -- 0x0221
        "00000010", -- 0x0222
        "00000011", -- 0x0223
        "00101000", -- 0x0224
        "10010000", -- 0x0225
        "00000001", -- 0x0226
        "01000100", -- 0x0227
        "11101001", -- 0x0228
        "11110000", -- 0x0229
        "10000000", -- 0x022A
        "10101101", -- 0x022B
        "01111000", -- 0x022C
        "00000000", -- 0x022D
        "10010000", -- 0x022E
        "00000001", -- 0x022F
        "00011010", -- 0x0230
        "01110100", -- 0x0231
        "00000110", -- 0x0232
        "11110000", -- 0x0233
        "00000010", -- 0x0234
        "00000011", -- 0x0235
        "00101000", -- 0x0236
        "00010010", -- 0x0237
        "00011100", -- 0x0238
        "10101011", -- 0x0239
        "10010000", -- 0x023A
        "00000001", -- 0x023B
        "00011010", -- 0x023C
        "01110100", -- 0x023D
        "00001001", -- 0x023E
        "11110000", -- 0x023F
        "00010010", -- 0x0240
        "00011001", -- 0x0241
        "01001000", -- 0x0242
        "10010000", -- 0x0243
        "00010111", -- 0x0244
        "11010011", -- 0x0245
        "00010010", -- 0x0246
        "00011101", -- 0x0247
        "00010001", -- 0x0248
        "10010000", -- 0x0249
        "00000001", -- 0x024A
        "00101101", -- 0x024B
        "00010010", -- 0x024C
        "00100001", -- 0x024D
        "11001000", -- 0x024E
        "10000000", -- 0x024F
        "10001000", -- 0x0250
        "00010010", -- 0x0251
        "00011101", -- 0x0252
        "10001011", -- 0x0253
        "11000100", -- 0x0254
        "00010010", -- 0x0255
        "00100000", -- 0x0256
        "00111001", -- 0x0257
        "00010010", -- 0x0258
        "00100001", -- 0x0259
        "00010001", -- 0x025A
        "00010010", -- 0x025B
        "00100001", -- 0x025C
        "01101000", -- 0x025D
        "11000011", -- 0x025E
        "00010011", -- 0x025F
        "01010100", -- 0x0260
        "01111100", -- 0x0261
        "10010000", -- 0x0262
        "00000001", -- 0x0263
        "01011010", -- 0x0264
        "11110000", -- 0x0265
        "00010010", -- 0x0266
        "00100100", -- 0x0267
        "01001000", -- 0x0268
        "00010010", -- 0x0269
        "00100100", -- 0x026A
        "01111000", -- 0x026B
        "11101111", -- 0x026C
        "00100101", -- 0x026D
        "11100000", -- 0x026E
        "10010000", -- 0x026F
        "00000001", -- 0x0270
        "01011011", -- 0x0271
        "00010010", -- 0x0272
        "00011100", -- 0x0273
        "11101111", -- 0x0274
        "00000010", -- 0x0275
        "00000001", -- 0x0276
        "11011001", -- 0x0277
        "00010010", -- 0x0278
        "00011101", -- 0x0279
        "10001011", -- 0x027A
        "00010010", -- 0x027B
        "00100000", -- 0x027C
        "00111001", -- 0x027D
        "11000100", -- 0x027E
        "00010010", -- 0x027F
        "00100001", -- 0x0280
        "00010001", -- 0x0281
        "11110000", -- 0x0282
        "10010000", -- 0x0283
        "00000001", -- 0x0284
        "01011010", -- 0x0285
        "11100100", -- 0x0286
        "00010010", -- 0x0287
        "00100001", -- 0x0288
        "01101000", -- 0x0289
        "00010010", -- 0x028A
        "00100100", -- 0x028B
        "01111000", -- 0x028C
        "10010000", -- 0x028D
        "00000001", -- 0x028E
        "01011011", -- 0x028F
        "11101111", -- 0x0290
        "00010010", -- 0x0291
        "00011100", -- 0x0292
        "11101111", -- 0x0293
        "00000010", -- 0x0294
        "00000001", -- 0x0295
        "11011001", -- 0x0296
        "11100100", -- 0x0297
        "11111101", -- 0x0298
        "11111100", -- 0x0299
        "01111110", -- 0x029A
        "00000100", -- 0x029B
        "01111111", -- 0x029C
        "11001101", -- 0x029D
        "00010010", -- 0x029E
        "00010100", -- 0x029F
        "00010100", -- 0x02A0
        "00010010", -- 0x02A1
        "00100010", -- 0x02A2
        "10101100", -- 0x02A3
        "01110101", -- 0x02A4
        "10110000", -- 0x02A5
        "00000000", -- 0x02A6
        "00000010", -- 0x02A7
        "00000001", -- 0x02A8
        "11011001", -- 0x02A9
        "01110101", -- 0x02AA
        "11100101", -- 0x02AB
        "11111111", -- 0x02AC
        "10000101", -- 0x02AD
        "00001100", -- 0x02AE
        "10000010", -- 0x02AF
        "10000101", -- 0x02B0
        "00001011", -- 0x02B1
        "10000011", -- 0x02B2
        "11100000", -- 0x02B3
        "01100100", -- 0x02B4
        "00010101", -- 0x02B5
        "01100000", -- 0x02B6
        "00000101", -- 0x02B7
        "01111111", -- 0x02B8
        "00000000", -- 0x02B9
        "00010010", -- 0x02BA
        "00011000", -- 0x02BB
        "01010010", -- 0x02BC
        "11100100", -- 0x02BD
        "11111110", -- 0x02BE
        "11111101", -- 0x02BF
        "11111100", -- 0x02C0
        "01111111", -- 0x02C1
        "01100100", -- 0x02C2
        "00010010", -- 0x02C3
        "00010110", -- 0x02C4
        "00110100", -- 0x02C5
        "00010010", -- 0x02C6
        "00100001", -- 0x02C7
        "11110110", -- 0x02C8
        "11110101", -- 0x02C9
        "11100101", -- 0x02CA
        "01111000", -- 0x02CB
        "11111111", -- 0x02CC
        "10000000", -- 0x02CD
        "01011001", -- 0x02CE
        "00010010", -- 0x02CF
        "00100001", -- 0x02D0
        "11110110", -- 0x02D1
        "11110101", -- 0x02D2
        "10110000", -- 0x02D3
        "00000010", -- 0x02D4
        "00000001", -- 0x02D5
        "11011001", -- 0x02D6
        "01010011", -- 0x02D7
        "11010101", -- 0x02D8
        "11110011", -- 0x02D9
        "01000011", -- 0x02DA
        "11010101", -- 0x02DB
        "00000100", -- 0x02DC
        "01010011", -- 0x02DD
        "11010101", -- 0x02DE
        "11001111", -- 0x02DF
        "01000011", -- 0x02E0
        "11010101", -- 0x02E1
        "00010000", -- 0x02E2
        "00000010", -- 0x02E3
        "00000001", -- 0x02E4
        "11011001", -- 0x02E5
        "00010010", -- 0x02E6
        "00100001", -- 0x02E7
        "11100000", -- 0x02E8
        "00000010", -- 0x02E9
        "00000001", -- 0x02EA
        "11011001", -- 0x02EB
        "00010010", -- 0x02EC
        "00100010", -- 0x02ED
        "10100011", -- 0x02EE
        "11100100", -- 0x02EF
        "11111101", -- 0x02F0
        "11111100", -- 0x02F1
        "01111110", -- 0x02F2
        "00011010", -- 0x02F3
        "01111111", -- 0x02F4
        "00101011", -- 0x02F5
        "00010010", -- 0x02F6
        "00010100", -- 0x02F7
        "00010100", -- 0x02F8
        "00000010", -- 0x02F9
        "00000001", -- 0x02FA
        "11011001", -- 0x02FB
        "00010010", -- 0x02FC
        "00011100", -- 0x02FD
        "10101011", -- 0x02FE
        "10010000", -- 0x02FF
        "00010111", -- 0x0300
        "11010101", -- 0x0301
        "11100000", -- 0x0302
        "11111100", -- 0x0303
        "10100011", -- 0x0304
        "11100000", -- 0x0305
        "11111101", -- 0x0306
        "01111110", -- 0x0307
        "00011010", -- 0x0308
        "01111111", -- 0x0309
        "00101011", -- 0x030A
        "00010010", -- 0x030B
        "00010100", -- 0x030C
        "00010100", -- 0x030D
        "00000010", -- 0x030E
        "00000001", -- 0x030F
        "11011001", -- 0x0310
        "00010010", -- 0x0311
        "00100001", -- 0x0312
        "11110110", -- 0x0313
        "11111000", -- 0x0314
        "01100000", -- 0x0315
        "00000100", -- 0x0316
        "10001000", -- 0x0317
        "00000001", -- 0x0318
        "11011001", -- 0x0319
        "00001011", -- 0x031A
        "10010000", -- 0x031B
        "00000001", -- 0x031C
        "01000010", -- 0x031D
        "11101000", -- 0x031E
        "11110000", -- 0x031F
        "00010010", -- 0x0320
        "00000011", -- 0x0321
        "00101010", -- 0x0322
        "00000010", -- 0x0323
        "00000001", -- 0x0324
        "11011001", -- 0x0325
        "01111000", -- 0x0326
        "11001100", -- 0x0327
        "11101000", -- 0x0328
        "00100010", -- 0x0329
        "11100101", -- 0x032A
        "11101101", -- 0x032B
        "00010010", -- 0x032C
        "00100010", -- 0x032D
        "01011110", -- 0x032E
        "01110000", -- 0x032F
        "00111100", -- 0x0330
        "00010010", -- 0x0331
        "00100011", -- 0x0332
        "01010110", -- 0x0333
        "01111111", -- 0x0334
        "00000011", -- 0x0335
        "00010010", -- 0x0336
        "00010001", -- 0x0337
        "11110101", -- 0x0338
        "00010010", -- 0x0339
        "00011001", -- 0x033A
        "01001000", -- 0x033B
        "10010000", -- 0x033C
        "00000001", -- 0x033D
        "00100101", -- 0x033E
        "00010010", -- 0x033F
        "00100001", -- 0x0340
        "11001000", -- 0x0341
        "10010000", -- 0x0342
        "00000001", -- 0x0343
        "10010011", -- 0x0344
        "00010010", -- 0x0345
        "00100100", -- 0x0346
        "01110011", -- 0x0347
        "10010000", -- 0x0348
        "00000001", -- 0x0349
        "00100001", -- 0x034A
        "00010010", -- 0x034B
        "00100100", -- 0x034C
        "01010100", -- 0x034D
        "10010000", -- 0x034E
        "00000001", -- 0x034F
        "10010110", -- 0x0350
        "11100000", -- 0x0351
        "10010000", -- 0x0352
        "00000000", -- 0x0353
        "00000101", -- 0x0354
        "11110000", -- 0x0355
        "10010000", -- 0x0356
        "00000001", -- 0x0357
        "00011111", -- 0x0358
        "00010010", -- 0x0359
        "00100100", -- 0x035A
        "01010100", -- 0x035B
        "01010011", -- 0x035C
        "11101101", -- 0x035D
        "11001111", -- 0x035E
        "10010000", -- 0x035F
        "00000001", -- 0x0360
        "01000010", -- 0x0361
        "11100000", -- 0x0362
        "00010010", -- 0x0363
        "00011110", -- 0x0364
        "00101101", -- 0x0365
        "01111100", -- 0x0366
        "00000000", -- 0x0367
        "01111101", -- 0x0368
        "01100100", -- 0x0369
        "00010010", -- 0x036A
        "00100011", -- 0x036B
        "01011110", -- 0x036C
        "10010000", -- 0x036D
        "00000001", -- 0x036E
        "00101001", -- 0x036F
        "11100100", -- 0x0370
        "11111111", -- 0x0371
        "11111110", -- 0x0372
        "11111101", -- 0x0373
        "11111100", -- 0x0374
        "00010010", -- 0x0375
        "00100001", -- 0x0376
        "11001000", -- 0x0377
        "10010000", -- 0x0378
        "00000001", -- 0x0379
        "01000000", -- 0x037A
        "00010010", -- 0x037B
        "00000000", -- 0x037C
        "00010110", -- 0x037D
        "01100000", -- 0x037E
        "00011111", -- 0x037F
        "00010010", -- 0x0380
        "00100010", -- 0x0381
        "11111101", -- 0x0382
        "10010000", -- 0x0383
        "00000001", -- 0x0384
        "00100001", -- 0x0385
        "11100000", -- 0x0386
        "11111100", -- 0x0387
        "10100011", -- 0x0388
        "11100000", -- 0x0389
        "11111101", -- 0x038A
        "00101001", -- 0x038B
        "11111001", -- 0x038C
        "11101000", -- 0x038D
        "00111100", -- 0x038E
        "11111000", -- 0x038F
        "11101011", -- 0x0390
        "11000011", -- 0x0391
        "10011001", -- 0x0392
        "11101010", -- 0x0393
        "10011000", -- 0x0394
        "01000000", -- 0x0395
        "00001000", -- 0x0396
        "00010010", -- 0x0397
        "00100011", -- 0x0398
        "00101110", -- 0x0399
        "01111111", -- 0x039A
        "00000001", -- 0x039B
        "00010010", -- 0x039C
        "00100001", -- 0x039D
        "11001000", -- 0x039E
        "00010010", -- 0x039F
        "00100010", -- 0x03A0
        "11111101", -- 0x03A1
        "10010000", -- 0x03A2
        "00000001", -- 0x03A3
        "01000011", -- 0x03A4
        "11100000", -- 0x03A5
        "11111000", -- 0x03A6
        "10010000", -- 0x03A7
        "00000001", -- 0x03A8
        "10001111", -- 0x03A9
        "11100000", -- 0x03AA
        "11010011", -- 0x03AB
        "10011000", -- 0x03AC
        "01000000", -- 0x03AD
        "00001000", -- 0x03AE
        "00010010", -- 0x03AF
        "00100011", -- 0x03B0
        "00101110", -- 0x03B1
        "01111111", -- 0x03B2
        "00000100", -- 0x03B3
        "00010010", -- 0x03B4
        "00100001", -- 0x03B5
        "11001000", -- 0x03B6
        "10010000", -- 0x03B7
        "00000001", -- 0x03B8
        "01000100", -- 0x03B9
        "11100000", -- 0x03BA
        "10110100", -- 0x03BB
        "00000001", -- 0x03BC
        "00011100", -- 0x03BD
        "11100101", -- 0x03BE
        "11011100", -- 0x03BF
        "00010010", -- 0x03C0
        "00100010", -- 0x03C1
        "01011110", -- 0x03C2
        "01110000", -- 0x03C3
        "00010101", -- 0x03C4
        "11100101", -- 0x03C5
        "11011100", -- 0x03C6
        "01010100", -- 0x03C7
        "00110000", -- 0x03C8
        "01100100", -- 0x03C9
        "00010000", -- 0x03CA
        "00100100", -- 0x03CB
        "11111111", -- 0x03CC
        "10110011", -- 0x03CD
        "11100100", -- 0x03CE
        "00110011", -- 0x03CF
        "01110000", -- 0x03D0
        "00001000", -- 0x03D1
        "00010010", -- 0x03D2
        "00100011", -- 0x03D3
        "00101110", -- 0x03D4
        "01111111", -- 0x03D5
        "00000101", -- 0x03D6
        "00010010", -- 0x03D7
        "00100001", -- 0x03D8
        "11001000", -- 0x03D9
        "10010000", -- 0x03DA
        "00000001", -- 0x03DB
        "00011111", -- 0x03DC
        "00010010", -- 0x03DD
        "00100100", -- 0x03DE
        "01110011", -- 0x03DF
        "11101011", -- 0x03E0
        "11010011", -- 0x03E1
        "10011001", -- 0x03E2
        "11101010", -- 0x03E3
        "10011000", -- 0x03E4
        "01000000", -- 0x03E5
        "01110100", -- 0x03E6
        "10010000", -- 0x03E7
        "00000001", -- 0x03E8
        "10010110", -- 0x03E9
        "11100000", -- 0x03EA
        "11111001", -- 0x03EB
        "11111111", -- 0x03EC
        "01111110", -- 0x03ED
        "00000000", -- 0x03EE
        "10010000", -- 0x03EF
        "00000000", -- 0x03F0
        "00000101", -- 0x03F1
        "11100000", -- 0x03F2
        "01111000", -- 0x03F3
        "00000000", -- 0x03F4
        "00100100", -- 0x03F5
        "00010100", -- 0x03F6
        "11111101", -- 0x03F7
        "11100100", -- 0x03F8
        "00111000", -- 0x03F9
        "11111100", -- 0x03FA
        "11101111", -- 0x03FB
        "11010011", -- 0x03FC
        "10011101", -- 0x03FD
        "11101110", -- 0x03FE
        "10011100", -- 0x03FF
        "00110000", -- 0x0400
        "11010010", -- 0x0401
        "00000010", -- 0x0402
        "10110010", -- 0x0403
        "11100111", -- 0x0404
        "00110000", -- 0x0405
        "11100111", -- 0x0406
        "01001110", -- 0x0407
        "10010000", -- 0x0408
        "00000001", -- 0x0409
        "00111101", -- 0x040A
        "11100000", -- 0x040B
        "11111000", -- 0x040C
        "01100000", -- 0x040D
        "01000111", -- 0x040E
        "10010000", -- 0x040F
        "00000001", -- 0x0410
        "01000101", -- 0x0411
        "11100000", -- 0x0412
        "00101000", -- 0x0413
        "11111101", -- 0x0414
        "11100100", -- 0x0415
        "00110011", -- 0x0416
        "11111100", -- 0x0417
        "11101101", -- 0x0418
        "11010011", -- 0x0419
        "10011111", -- 0x041A
        "11101100", -- 0x041B
        "10011110", -- 0x041C
        "00110000", -- 0x041D
        "11010010", -- 0x041E
        "00000010", -- 0x041F
        "10110010", -- 0x0420
        "11100111", -- 0x0421
        "00110000", -- 0x0422
        "11100111", -- 0x0423
        "00110001", -- 0x0424
        "11101001", -- 0x0425
        "00010010", -- 0x0426
        "00100100", -- 0x0427
        "01000010", -- 0x0428
        "10010000", -- 0x0429
        "00010111", -- 0x042A
        "11010111", -- 0x042B
        "00010010", -- 0x042C
        "00100001", -- 0x042D
        "11001000", -- 0x042E
        "11101001", -- 0x042F
        "00010010", -- 0x0430
        "00100100", -- 0x0431
        "01000010", -- 0x0432
        "01110100", -- 0x0433
        "00010000", -- 0x0434
        "00010010", -- 0x0435
        "00011111", -- 0x0436
        "00110000", -- 0x0437
        "10010000", -- 0x0438
        "00010111", -- 0x0439
        "11010111", -- 0x043A
        "00010010", -- 0x043B
        "00100001", -- 0x043C
        "11001000", -- 0x043D
        "11100100", -- 0x043E
        "11111110", -- 0x043F
        "11111101", -- 0x0440
        "11111100", -- 0x0441
        "10010000", -- 0x0442
        "00010111", -- 0x0443
        "11010111", -- 0x0444
        "01111111", -- 0x0445
        "00000011", -- 0x0446
        "00010010", -- 0x0447
        "00011011", -- 0x0448
        "11010001", -- 0x0449
        "10010000", -- 0x044A
        "00010111", -- 0x044B
        "11010111", -- 0x044C
        "00010010", -- 0x044D
        "00100001", -- 0x044E
        "10111100", -- 0x044F
        "10010000", -- 0x0450
        "00000001", -- 0x0451
        "00101001", -- 0x0452
        "00010010", -- 0x0453
        "00100001", -- 0x0454
        "11001000", -- 0x0455
        "10010000", -- 0x0456
        "00000000", -- 0x0457
        "00000101", -- 0x0458
        "11101001", -- 0x0459
        "11110000", -- 0x045A
        "10010000", -- 0x045B
        "00000001", -- 0x045C
        "00011111", -- 0x045D
        "11101010", -- 0x045E
        "11110000", -- 0x045F
        "11101011", -- 0x0460
        "10100011", -- 0x0461
        "11110000", -- 0x0462
        "10010000", -- 0x0463
        "00000001", -- 0x0464
        "00111110", -- 0x0465
        "00010010", -- 0x0466
        "00000000", -- 0x0467
        "00010110", -- 0x0468
        "01100000", -- 0x0469
        "00111000", -- 0x046A
        "00010010", -- 0x046B
        "00011001", -- 0x046C
        "01001000", -- 0x046D
        "10010000", -- 0x046E
        "00010111", -- 0x046F
        "11011011", -- 0x0470
        "00010010", -- 0x0471
        "00100001", -- 0x0472
        "11001000", -- 0x0473
        "10010000", -- 0x0474
        "00000001", -- 0x0475
        "00100101", -- 0x0476
        "00010010", -- 0x0477
        "00100001", -- 0x0478
        "10111100", -- 0x0479
        "10010000", -- 0x047A
        "00010111", -- 0x047B
        "11011011", -- 0x047C
        "00010010", -- 0x047D
        "00011011", -- 0x047E
        "01011101", -- 0x047F
        "11100100", -- 0x0480
        "11111101", -- 0x0481
        "11111100", -- 0x0482
        "10010000", -- 0x0483
        "00010111", -- 0x0484
        "11011011", -- 0x0485
        "01111110", -- 0x0486
        "00000011", -- 0x0487
        "01111111", -- 0x0488
        "11101000", -- 0x0489
        "00010010", -- 0x048A
        "00011010", -- 0x048B
        "01011110", -- 0x048C
        "10010000", -- 0x048D
        "00000001", -- 0x048E
        "00111110", -- 0x048F
        "00010010", -- 0x0490
        "00100011", -- 0x0491
        "01000110", -- 0x0492
        "10010000", -- 0x0493
        "00010111", -- 0x0494
        "11011011", -- 0x0495
        "00010010", -- 0x0496
        "00100011", -- 0x0497
        "10100100", -- 0x0498
        "01000000", -- 0x0499
        "00001000", -- 0x049A
        "00010010", -- 0x049B
        "00100011", -- 0x049C
        "00101110", -- 0x049D
        "01111111", -- 0x049E
        "00000010", -- 0x049F
        "00010010", -- 0x04A0
        "00100001", -- 0x04A1
        "11001000", -- 0x04A2
        "11100100", -- 0x04A3
        "11111111", -- 0x04A4
        "11111110", -- 0x04A5
        "11111101", -- 0x04A6
        "11111100", -- 0x04A7
        "10010000", -- 0x04A8
        "00000001", -- 0x04A9
        "00101001", -- 0x04AA
        "00010010", -- 0x04AB
        "00100011", -- 0x04AC
        "10100100", -- 0x04AD
        "01100000", -- 0x04AE
        "00011100", -- 0x04AF
        "01000000", -- 0x04B0
        "00011010", -- 0x04B1
        "11100100", -- 0x04B2
        "11111101", -- 0x04B3
        "11111100", -- 0x04B4
        "00010010", -- 0x04B5
        "00100011", -- 0x04B6
        "01011110", -- 0x04B7
        "00010010", -- 0x04B8
        "00100011", -- 0x04B9
        "11000111", -- 0x04BA
        "10010000", -- 0x04BB
        "00000001", -- 0x04BC
        "00101001", -- 0x04BD
        "00010010", -- 0x04BE
        "00100001", -- 0x04BF
        "10111100", -- 0x04C0
        "00010010", -- 0x04C1
        "00100100", -- 0x04C2
        "00010010", -- 0x04C3
        "01111111", -- 0x04C4
        "00000100", -- 0x04C5
        "00010010", -- 0x04C6
        "00010001", -- 0x04C7
        "11110101", -- 0x04C8
        "00010010", -- 0x04C9
        "00100010", -- 0x04CA
        "10100011", -- 0x04CB
        "00100010", -- 0x04CC
        "00010010", -- 0x04CD
        "00100100", -- 0x04CE
        "00001100", -- 0x04CF
        "01001000", -- 0x04D0
        "01110000", -- 0x04D1
        "00011111", -- 0x04D2
        "00010010", -- 0x04D3
        "00100010", -- 0x04D4
        "00100010", -- 0x04D5
        "11100100", -- 0x04D6
        "11110000", -- 0x04D7
        "10100011", -- 0x04D8
        "11110000", -- 0x04D9
        "10010000", -- 0x04DA
        "00000001", -- 0x04DB
        "01011100", -- 0x04DC
        "01110100", -- 0x04DD
        "00000001", -- 0x04DE
        "11110000", -- 0x04DF
        "01110101", -- 0x04E0
        "10110000", -- 0x04E1
        "00000000", -- 0x04E2
        "10010000", -- 0x04E3
        "00000001", -- 0x04E4
        "01010001", -- 0x04E5
        "11100000", -- 0x04E6
        "00010010", -- 0x04E7
        "00100100", -- 0x04E8
        "01000010", -- 0x04E9
        "00010010", -- 0x04EA
        "00100100", -- 0x04EB
        "00010010", -- 0x04EC
        "01111111", -- 0x04ED
        "00001011", -- 0x04EE
        "00010010", -- 0x04EF
        "00010001", -- 0x04F0
        "11110101", -- 0x04F1
        "01010011", -- 0x04F2
        "11010101", -- 0x04F3
        "11001111", -- 0x04F4
        "01000011", -- 0x04F5
        "11010101", -- 0x04F6
        "00010000", -- 0x04F7
        "01110101", -- 0x04F8
        "11010100", -- 0x04F9
        "00000001", -- 0x04FA
        "00010010", -- 0x04FB
        "00100000", -- 0x04FC
        "01011001", -- 0x04FD
        "10010000", -- 0x04FE
        "00000001", -- 0x04FF
        "10101111", -- 0x0500
        "00010010", -- 0x0501
        "00100100", -- 0x0502
        "01010100", -- 0x0503
        "10010000", -- 0x0504
        "00000001", -- 0x0505
        "10101111", -- 0x0506
        "00010010", -- 0x0507
        "00100010", -- 0x0508
        "10110101", -- 0x0509
        "10010000", -- 0x050A
        "00000001", -- 0x050B
        "10101111", -- 0x050C
        "01111110", -- 0x050D
        "00000000", -- 0x050E
        "00010010", -- 0x050F
        "00011111", -- 0x0510
        "10010001", -- 0x0511
        "01010011", -- 0x0512
        "11010101", -- 0x0513
        "11001111", -- 0x0514
        "01000011", -- 0x0515
        "11010101", -- 0x0516
        "00100000", -- 0x0517
        "01010011", -- 0x0518
        "11010101", -- 0x0519
        "11110011", -- 0x051A
        "01000011", -- 0x051B
        "11010101", -- 0x051C
        "00000100", -- 0x051D
        "01110101", -- 0x051E
        "11010100", -- 0x051F
        "00000011", -- 0x0520
        "00010010", -- 0x0521
        "00100000", -- 0x0522
        "01011001", -- 0x0523
        "10010000", -- 0x0524
        "00000001", -- 0x0525
        "10101101", -- 0x0526
        "00010010", -- 0x0527
        "00100100", -- 0x0528
        "01010100", -- 0x0529
        "10010000", -- 0x052A
        "00000001", -- 0x052B
        "10101101", -- 0x052C
        "00010010", -- 0x052D
        "00100010", -- 0x052E
        "10110101", -- 0x052F
        "10010000", -- 0x0530
        "00000001", -- 0x0531
        "10101101", -- 0x0532
        "01111110", -- 0x0533
        "00000000", -- 0x0534
        "00010010", -- 0x0535
        "00011111", -- 0x0536
        "10010001", -- 0x0537
        "01010011", -- 0x0538
        "11010101", -- 0x0539
        "11110011", -- 0x053A
        "01000011", -- 0x053B
        "11010101", -- 0x053C
        "00001000", -- 0x053D
        "01110101", -- 0x053E
        "11010100", -- 0x053F
        "00000000", -- 0x0540
        "10010000", -- 0x0541
        "00000001", -- 0x0542
        "10101101", -- 0x0543
        "11100000", -- 0x0544
        "11111110", -- 0x0545
        "10100011", -- 0x0546
        "11100000", -- 0x0547
        "11111111", -- 0x0548
        "10100011", -- 0x0549
        "11100000", -- 0x054A
        "11111100", -- 0x054B
        "10100011", -- 0x054C
        "11100000", -- 0x054D
        "11111101", -- 0x054E
        "00010010", -- 0x054F
        "00010011", -- 0x0550
        "01000100", -- 0x0551
        "10010000", -- 0x0552
        "00000001", -- 0x0553
        "01010001", -- 0x0554
        "11100000", -- 0x0555
        "10110100", -- 0x0556
        "00001100", -- 0x0557
        "00000010", -- 0x0558
        "10000000", -- 0x0559
        "00000011", -- 0x055A
        "00000010", -- 0x055B
        "00000110", -- 0x055C
        "00011110", -- 0x055D
        "10010000", -- 0x055E
        "00000001", -- 0x055F
        "01010100", -- 0x0560
        "00010010", -- 0x0561
        "00000000", -- 0x0562
        "00010110", -- 0x0563
        "01110000", -- 0x0564
        "00000011", -- 0x0565
        "00000010", -- 0x0566
        "00000101", -- 0x0567
        "11111110", -- 0x0568
        "10010000", -- 0x0569
        "00000001", -- 0x056A
        "01011100", -- 0x056B
        "11100000", -- 0x056C
        "01111000", -- 0x056D
        "00000000", -- 0x056E
        "01010100", -- 0x056F
        "00000001", -- 0x0570
        "11111011", -- 0x0571
        "11100100", -- 0x0572
        "11111010", -- 0x0573
        "01001011", -- 0x0574
        "01100000", -- 0x0575
        "00011011", -- 0x0576
        "11100101", -- 0x0577
        "10110000", -- 0x0578
        "01110000", -- 0x0579
        "00001111", -- 0x057A
        "10010000", -- 0x057B
        "00000001", -- 0x057C
        "01011010", -- 0x057D
        "11100000", -- 0x057E
        "00010010", -- 0x057F
        "00100100", -- 0x0580
        "01000010", -- 0x0581
        "00010010", -- 0x0582
        "00100100", -- 0x0583
        "00010010", -- 0x0584
        "01111111", -- 0x0585
        "00001111", -- 0x0586
        "00010010", -- 0x0587
        "00010001", -- 0x0588
        "11110101", -- 0x0589
        "10010000", -- 0x058A
        "00000001", -- 0x058B
        "01011010", -- 0x058C
        "11100000", -- 0x058D
        "11110101", -- 0x058E
        "10110000", -- 0x058F
        "10000000", -- 0x0590
        "00010000", -- 0x0591
        "10101000", -- 0x0592
        "10110000", -- 0x0593
        "11101000", -- 0x0594
        "01100000", -- 0x0595
        "00001000", -- 0x0596
        "00010010", -- 0x0597
        "00100011", -- 0x0598
        "01010110", -- 0x0599
        "01111111", -- 0x059A
        "00010000", -- 0x059B
        "00010010", -- 0x059C
        "00010001", -- 0x059D
        "11110101", -- 0x059E
        "01110101", -- 0x059F
        "10110000", -- 0x05A0
        "00000000", -- 0x05A1
        "00010010", -- 0x05A2
        "00100100", -- 0x05A3
        "00001100", -- 0x05A4
        "11111001", -- 0x05A5
        "10010000", -- 0x05A6
        "00000001", -- 0x05A7
        "01010110", -- 0x05A8
        "00010010", -- 0x05A9
        "00100010", -- 0x05AA
        "00001100", -- 0x05AB
        "01000000", -- 0x05AC
        "01000000", -- 0x05AD
        "00010010", -- 0x05AE
        "00100001", -- 0x05AF
        "01000100", -- 0x05B0
        "01000000", -- 0x05B1
        "00011100", -- 0x05B2
        "10010000", -- 0x05B3
        "00000001", -- 0x05B4
        "01011011", -- 0x05B5
        "00010010", -- 0x05B6
        "00100100", -- 0x05B7
        "10000111", -- 0x05B8
        "11000011", -- 0x05B9
        "10011000", -- 0x05BA
        "01000000", -- 0x05BB
        "00001001", -- 0x05BC
        "00010010", -- 0x05BD
        "00100100", -- 0x05BE
        "01001110", -- 0x05BF
        "01110101", -- 0x05C0
        "10110000", -- 0x05C1
        "00000000", -- 0x05C2
        "00000010", -- 0x05C3
        "00011111", -- 0x05C4
        "10100011", -- 0x05C5
        "00010010", -- 0x05C6
        "00100011", -- 0x05C7
        "11111000", -- 0x05C8
        "00010010", -- 0x05C9
        "00100010", -- 0x05CA
        "00101100", -- 0x05CB
        "00000010", -- 0x05CC
        "00011110", -- 0x05CD
        "11001011", -- 0x05CE
        "00010010", -- 0x05CF
        "00100010", -- 0x05D0
        "00100010", -- 0x05D1
        "00010010", -- 0x05D2
        "00011111", -- 0x05D3
        "01011000", -- 0x05D4
        "00010010", -- 0x05D5
        "00100001", -- 0x05D6
        "00101011", -- 0x05D7
        "10001111", -- 0x05D8
        "00011011", -- 0x05D9
        "10001110", -- 0x05DA
        "00011010", -- 0x05DB
        "00010010", -- 0x05DC
        "00100011", -- 0x05DD
        "11111111", -- 0x05DE
        "10101111", -- 0x05DF
        "00011011", -- 0x05E0
        "10101110", -- 0x05E1
        "00011010", -- 0x05E2
        "00010010", -- 0x05E3
        "00100100", -- 0x05E4
        "10010101", -- 0x05E5
        "00010010", -- 0x05E6
        "00100100", -- 0x05E7
        "00010010", -- 0x05E8
        "01111111", -- 0x05E9
        "00001101", -- 0x05EA
        "00000010", -- 0x05EB
        "00010001", -- 0x05EC
        "11110101", -- 0x05ED
        "00010010", -- 0x05EE
        "00100001", -- 0x05EF
        "00101011", -- 0x05F0
        "10001111", -- 0x05F1
        "00000101", -- 0x05F2
        "10001110", -- 0x05F3
        "00000100", -- 0x05F4
        "10010000", -- 0x05F5
        "00000001", -- 0x05F6
        "01011000", -- 0x05F7
        "00010010", -- 0x05F8
        "00011111", -- 0x05F9
        "01011000", -- 0x05FA
        "00000010", -- 0x05FB
        "00100011", -- 0x05FC
        "01101100", -- 0x05FD
        "00010010", -- 0x05FE
        "00100100", -- 0x05FF
        "00001100", -- 0x0600
        "00100100", -- 0x0601
        "11110000", -- 0x0602
        "11101000", -- 0x0603
        "00110100", -- 0x0604
        "11111111", -- 0x0605
        "01010000", -- 0x0606
        "00001001", -- 0x0607
        "00010010", -- 0x0608
        "00100010", -- 0x0609
        "00101100", -- 0x060A
        "00010010", -- 0x060B
        "00100011", -- 0x060C
        "11010101", -- 0x060D
        "00000010", -- 0x060E
        "00100011", -- 0x060F
        "11111000", -- 0x0610
        "10010000", -- 0x0611
        "00000001", -- 0x0612
        "01011000", -- 0x0613
        "00010010", -- 0x0614
        "00011111", -- 0x0615
        "01011000", -- 0x0616
        "01111100", -- 0x0617
        "00000110", -- 0x0618
        "01111101", -- 0x0619
        "01000000", -- 0x061A
        "00000010", -- 0x061B
        "00100011", -- 0x061C
        "01101100", -- 0x061D
        "10010000", -- 0x061E
        "00000001", -- 0x061F
        "01010110", -- 0x0620
        "11100000", -- 0x0621
        "11111100", -- 0x0622
        "10100011", -- 0x0623
        "11100000", -- 0x0624
        "11111101", -- 0x0625
        "01111110", -- 0x0626
        "00000000", -- 0x0627
        "01111111", -- 0x0628
        "11001000", -- 0x0629
        "00010010", -- 0x062A
        "00011110", -- 0x062B
        "10110110", -- 0x062C
        "00010010", -- 0x062D
        "00100011", -- 0x062E
        "11111111", -- 0x062F
        "10010000", -- 0x0630
        "00000001", -- 0x0631
        "01010100", -- 0x0632
        "00010010", -- 0x0633
        "00100100", -- 0x0634
        "10000111", -- 0x0635
        "01001000", -- 0x0636
        "01110000", -- 0x0637
        "00000110", -- 0x0638
        "10010000", -- 0x0639
        "00000001", -- 0x063A
        "01010100", -- 0x063B
        "00010010", -- 0x063C
        "00100011", -- 0x063D
        "11010101", -- 0x063E
        "00010010", -- 0x063F
        "00100001", -- 0x0640
        "01000100", -- 0x0641
        "01000000", -- 0x0642
        "00010101", -- 0x0643
        "10010000", -- 0x0644
        "00000001", -- 0x0645
        "01011011", -- 0x0646
        "00010010", -- 0x0647
        "00100100", -- 0x0648
        "10000111", -- 0x0649
        "10110101", -- 0x064A
        "00000000", -- 0x064B
        "00000110", -- 0x064C
        "00010010", -- 0x064D
        "00100100", -- 0x064E
        "01001110", -- 0x064F
        "00000010", -- 0x0650
        "00011111", -- 0x0651
        "10100011", -- 0x0652
        "10010000", -- 0x0653
        "00000001", -- 0x0654
        "01010100", -- 0x0655
        "00000010", -- 0x0656
        "00011110", -- 0x0657
        "11001011", -- 0x0658
        "10010000", -- 0x0659
        "00000001", -- 0x065A
        "01010100", -- 0x065B
        "00000010", -- 0x065C
        "00011111", -- 0x065D
        "01011000", -- 0x065E
        "00100010", -- 0x065F
        "10010000", -- 0x0660
        "00011111", -- 0x0661
        "11101000", -- 0x0662
        "11100100", -- 0x0663
        "10010011", -- 0x0664
        "01100000", -- 0x0665
        "11111000", -- 0x0666
        "11111111", -- 0x0667
        "10100011", -- 0x0668
        "11100100", -- 0x0669
        "10010011", -- 0x066A
        "10100011", -- 0x066B
        "11111110", -- 0x066C
        "11100100", -- 0x066D
        "10010011", -- 0x066E
        "10100011", -- 0x066F
        "11111000", -- 0x0670
        "11100100", -- 0x0671
        "10010011", -- 0x0672
        "10100011", -- 0x0673
        "11111001", -- 0x0674
        "11100100", -- 0x0675
        "10010011", -- 0x0676
        "10100011", -- 0x0677
        "11111010", -- 0x0678
        "11100100", -- 0x0679
        "10010011", -- 0x067A
        "10100011", -- 0x067B
        "11111011", -- 0x067C
        "11100100", -- 0x067D
        "10010011", -- 0x067E
        "10100011", -- 0x067F
        "11111100", -- 0x0680
        "11100100", -- 0x0681
        "10010011", -- 0x0682
        "11111101", -- 0x0683
        "10100011", -- 0x0684
        "11101110", -- 0x0685
        "01010100", -- 0x0686
        "00000001", -- 0x0687
        "01110000", -- 0x0688
        "01000110", -- 0x0689
        "11101111", -- 0x068A
        "01100100", -- 0x068B
        "00000001", -- 0x068C
        "01100000", -- 0x068D
        "00110011", -- 0x068E
        "11101111", -- 0x068F
        "01100100", -- 0x0690
        "00000011", -- 0x0691
        "01100000", -- 0x0692
        "00101110", -- 0x0693
        "10111111", -- 0x0694
        "00001001", -- 0x0695
        "00000010", -- 0x0696
        "10000000", -- 0x0697
        "00101001", -- 0x0698
        "10111111", -- 0x0699
        "00000100", -- 0x069A
        "00000111", -- 0x069B
        "10101110", -- 0x069C
        "10000011", -- 0x069D
        "10101111", -- 0x069E
        "10000010", -- 0x069F
        "00000010", -- 0x06A0
        "00000111", -- 0x06A1
        "01000110", -- 0x06A2
        "10111111", -- 0x06A3
        "00000110", -- 0x06A4
        "00000010", -- 0x06A5
        "10000000", -- 0x06A6
        "00100001", -- 0x06A7
        "10101110", -- 0x06A8
        "10000011", -- 0x06A9
        "10101111", -- 0x06AA
        "10000010", -- 0x06AB
        "10001000", -- 0x06AC
        "10000011", -- 0x06AD
        "10001001", -- 0x06AE
        "10000010", -- 0x06AF
        "11100100", -- 0x06B0
        "11110000", -- 0x06B1
        "10100011", -- 0x06B2
        "00011101", -- 0x06B3
        "10111101", -- 0x06B4
        "11111111", -- 0x06B5
        "00000001", -- 0x06B6
        "00011100", -- 0x06B7
        "11101100", -- 0x06B8
        "01001101", -- 0x06B9
        "01110000", -- 0x06BA
        "11110100", -- 0x06BB
        "10001110", -- 0x06BC
        "10000011", -- 0x06BD
        "10001111", -- 0x06BE
        "10000010", -- 0x06BF
        "10000000", -- 0x06C0
        "10100001", -- 0x06C1
        "11100100", -- 0x06C2
        "11110111", -- 0x06C3
        "00001001", -- 0x06C4
        "11011101", -- 0x06C5
        "11111011", -- 0x06C6
        "10000000", -- 0x06C7
        "10011010", -- 0x06C8
        "11100100", -- 0x06C9
        "11110011", -- 0x06CA
        "00001001", -- 0x06CB
        "11011101", -- 0x06CC
        "11111011", -- 0x06CD
        "10000000", -- 0x06CE
        "10010011", -- 0x06CF
        "11101111", -- 0x06D0
        "01100100", -- 0x06D1
        "00000001", -- 0x06D2
        "01100000", -- 0x06D3
        "01000101", -- 0x06D4
        "11101111", -- 0x06D5
        "01100100", -- 0x06D6
        "00000011", -- 0x06D7
        "01100000", -- 0x06D8
        "01000000", -- 0x06D9
        "10111111", -- 0x06DA
        "00001001", -- 0x06DB
        "00000010", -- 0x06DC
        "10000000", -- 0x06DD
        "00111011", -- 0x06DE
        "10111111", -- 0x06DF
        "00000100", -- 0x06E0
        "00001010", -- 0x06E1
        "10101110", -- 0x06E2
        "10000011", -- 0x06E3
        "10101111", -- 0x06E4
        "10000010", -- 0x06E5
        "10001010", -- 0x06E6
        "10000011", -- 0x06E7
        "10001011", -- 0x06E8
        "10000010", -- 0x06E9
        "10000000", -- 0x06EA
        "01011010", -- 0x06EB
        "10111111", -- 0x06EC
        "00000110", -- 0x06ED
        "00000010", -- 0x06EE
        "10000000", -- 0x06EF
        "00111111", -- 0x06F0
        "10101110", -- 0x06F1
        "10000011", -- 0x06F2
        "10101111", -- 0x06F3
        "10000010", -- 0x06F4
        "10001010", -- 0x06F5
        "10000011", -- 0x06F6
        "10001011", -- 0x06F7
        "10000010", -- 0x06F8
        "11100100", -- 0x06F9
        "10010011", -- 0x06FA
        "10100011", -- 0x06FB
        "10101010", -- 0x06FC
        "10000011", -- 0x06FD
        "10101011", -- 0x06FE
        "10000010", -- 0x06FF
        "10001000", -- 0x0700
        "10000011", -- 0x0701
        "10001001", -- 0x0702
        "10000010", -- 0x0703
        "11110000", -- 0x0704
        "10100011", -- 0x0705
        "10101000", -- 0x0706
        "10000011", -- 0x0707
        "10101001", -- 0x0708
        "10000010", -- 0x0709
        "00011101", -- 0x070A
        "10111101", -- 0x070B
        "11111111", -- 0x070C
        "00000001", -- 0x070D
        "00011100", -- 0x070E
        "11101100", -- 0x070F
        "01001101", -- 0x0710
        "01110000", -- 0x0711
        "11100010", -- 0x0712
        "10001110", -- 0x0713
        "10000011", -- 0x0714
        "10001111", -- 0x0715
        "10000010", -- 0x0716
        "00000010", -- 0x0717
        "00000110", -- 0x0718
        "01100011", -- 0x0719
        "10101110", -- 0x071A
        "10000011", -- 0x071B
        "10101111", -- 0x071C
        "10000010", -- 0x071D
        "10001010", -- 0x071E
        "10000011", -- 0x071F
        "10001011", -- 0x0720
        "10000010", -- 0x0721
        "11100100", -- 0x0722
        "10010011", -- 0x0723
        "11110111", -- 0x0724
        "00001001", -- 0x0725
        "10100011", -- 0x0726
        "11011101", -- 0x0727
        "11111001", -- 0x0728
        "10001110", -- 0x0729
        "10000011", -- 0x072A
        "10001111", -- 0x072B
        "10000010", -- 0x072C
        "00000010", -- 0x072D
        "00000110", -- 0x072E
        "01100011", -- 0x072F
        "10101110", -- 0x0730
        "10000011", -- 0x0731
        "10101111", -- 0x0732
        "10000010", -- 0x0733
        "10001010", -- 0x0734
        "10000011", -- 0x0735
        "10001011", -- 0x0736
        "10000010", -- 0x0737
        "11100100", -- 0x0738
        "10010011", -- 0x0739
        "11110011", -- 0x073A
        "00001001", -- 0x073B
        "10100011", -- 0x073C
        "11011101", -- 0x073D
        "11111001", -- 0x073E
        "10001110", -- 0x073F
        "10000011", -- 0x0740
        "10001111", -- 0x0741
        "10000010", -- 0x0742
        "00000010", -- 0x0743
        "00000110", -- 0x0744
        "01100011", -- 0x0745
        "11101001", -- 0x0746
        "01110101", -- 0x0747
        "11110000", -- 0x0748
        "00001000", -- 0x0749
        "10000100", -- 0x074A
        "00100100", -- 0x074B
        "00100000", -- 0x074C
        "11111000", -- 0x074D
        "11100110", -- 0x074E
        "11111100", -- 0x074F
        "11100101", -- 0x0750
        "11110000", -- 0x0751
        "01100000", -- 0x0752
        "00000101", -- 0x0753
        "11001100", -- 0x0754
        "00000011", -- 0x0755
        "11011100", -- 0x0756
        "11111101", -- 0x0757
        "11001100", -- 0x0758
        "10111101", -- 0x0759
        "00000000", -- 0x075A
        "00010100", -- 0x075B
        "11101001", -- 0x075C
        "01010100", -- 0x075D
        "00000111", -- 0x075E
        "01100000", -- 0x075F
        "00000110", -- 0x0760
        "11101100", -- 0x0761
        "00000011", -- 0x0762
        "11111100", -- 0x0763
        "00001001", -- 0x0764
        "10000000", -- 0x0765
        "11110101", -- 0x0766
        "11101100", -- 0x0767
        "11110110", -- 0x0768
        "10001110", -- 0x0769
        "10000011", -- 0x076A
        "10001111", -- 0x076B
        "10000010", -- 0x076C
        "00000010", -- 0x076D
        "00000110", -- 0x076E
        "01100011", -- 0x076F
        "11101011", -- 0x0770
        "01001010", -- 0x0771
        "01100000", -- 0x0772
        "00000011", -- 0x0773
        "11100100", -- 0x0774
        "10010011", -- 0x0775
        "10100011", -- 0x0776
        "11000011", -- 0x0777
        "01100000", -- 0x0778
        "00000001", -- 0x0779
        "11010011", -- 0x077A
        "11101100", -- 0x077B
        "00010011", -- 0x077C
        "11111100", -- 0x077D
        "00001001", -- 0x077E
        "00011101", -- 0x077F
        "11101001", -- 0x0780
        "01010100", -- 0x0781
        "00000111", -- 0x0782
        "01110000", -- 0x0783
        "11010100", -- 0x0784
        "11101100", -- 0x0785
        "11110110", -- 0x0786
        "10000000", -- 0x0787
        "10111101", -- 0x0788
        "00001111", -- 0x0789
        "10111111", -- 0x078A
        "00000000", -- 0x078B
        "00000001", -- 0x078C
        "00001110", -- 0x078D
        "10001111", -- 0x078E
        "00001100", -- 0x078F
        "10001110", -- 0x0790
        "00001011", -- 0x0791
        "10001111", -- 0x0792
        "10000010", -- 0x0793
        "10001110", -- 0x0794
        "10000011", -- 0x0795
        "11100000", -- 0x0796
        "00010010", -- 0x0797
        "00100100", -- 0x0798
        "01000010", -- 0x0799
        "00010010", -- 0x079A
        "00100100", -- 0x079B
        "00010010", -- 0x079C
        "01111111", -- 0x079D
        "00001010", -- 0x079E
        "00010010", -- 0x079F
        "00010001", -- 0x07A0
        "11110101", -- 0x07A1
        "10000101", -- 0x07A2
        "00001100", -- 0x07A3
        "10000010", -- 0x07A4
        "10000101", -- 0x07A5
        "00001011", -- 0x07A6
        "10000011", -- 0x07A7
        "11100000", -- 0x07A8
        "00010100", -- 0x07A9
        "01100000", -- 0x07AA
        "00010101", -- 0x07AB
        "00010100", -- 0x07AC
        "01110000", -- 0x07AD
        "00000011", -- 0x07AE
        "00000010", -- 0x07AF
        "00001000", -- 0x07B0
        "01000001", -- 0x07B1
        "00010100", -- 0x07B2
        "01100000", -- 0x07B3
        "01011111", -- 0x07B4
        "00010100", -- 0x07B5
        "01100000", -- 0x07B6
        "01101001", -- 0x07B7
        "00010100", -- 0x07B8
        "01110000", -- 0x07B9
        "00000011", -- 0x07BA
        "00000010", -- 0x07BB
        "00001000", -- 0x07BC
        "01101111", -- 0x07BD
        "00000010", -- 0x07BE
        "00001000", -- 0x07BF
        "10010011", -- 0x07C0
        "00010010", -- 0x07C1
        "00100011", -- 0x07C2
        "00011110", -- 0x07C3
        "00010010", -- 0x07C4
        "00100100", -- 0x07C5
        "01111101", -- 0x07C6
        "10010000", -- 0x07C7
        "00011000", -- 0x07C8
        "00001000", -- 0x07C9
        "01110100", -- 0x07CA
        "10100000", -- 0x07CB
        "11110000", -- 0x07CC
        "00010010", -- 0x07CD
        "00100011", -- 0x07CE
        "01111010", -- 0x07CF
        "01110100", -- 0x07D0
        "00010000", -- 0x07D1
        "00010010", -- 0x07D2
        "00100010", -- 0x07D3
        "00110110", -- 0x07D4
        "10100011", -- 0x07D5
        "01110100", -- 0x07D6
        "00101000", -- 0x07D7
        "00010010", -- 0x07D8
        "00100100", -- 0x07D9
        "01100100", -- 0x07DA
        "01110100", -- 0x07DB
        "10010110", -- 0x07DC
        "00010010", -- 0x07DD
        "00100100", -- 0x07DE
        "01011111", -- 0x07DF
        "00010100", -- 0x07E0
        "00010010", -- 0x07E1
        "00100100", -- 0x07E2
        "01011010", -- 0x07E3
        "10100011", -- 0x07E4
        "11100100", -- 0x07E5
        "00010010", -- 0x07E6
        "00100100", -- 0x07E7
        "01100100", -- 0x07E8
        "01110100", -- 0x07E9
        "00000010", -- 0x07EA
        "00010010", -- 0x07EB
        "00100010", -- 0x07EC
        "11010000", -- 0x07ED
        "00010010", -- 0x07EE
        "00100100", -- 0x07EF
        "00110000", -- 0x07F0
        "00010010", -- 0x07F1
        "00100100", -- 0x07F2
        "01011111", -- 0x07F3
        "00010010", -- 0x07F4
        "00100011", -- 0x07F5
        "00001110", -- 0x07F6
        "00010010", -- 0x07F7
        "00100100", -- 0x07F8
        "00110110", -- 0x07F9
        "00010010", -- 0x07FA
        "00100010", -- 0x07FB
        "00110110", -- 0x07FC
        "11100100", -- 0x07FD
        "11110000", -- 0x07FE
        "10100011", -- 0x07FF
        "01110100", -- 0x0800
        "00101000", -- 0x0801
        "00010010", -- 0x0802
        "00100010", -- 0x0803
        "11010000", -- 0x0804
        "01110100", -- 0x0805
        "00101010", -- 0x0806
        "11110000", -- 0x0807
        "10100011", -- 0x0808
        "01110100", -- 0x0809
        "00110000", -- 0x080A
        "00010010", -- 0x080B
        "00100011", -- 0x080C
        "00010110", -- 0x080D
        "00010010", -- 0x080E
        "00100100", -- 0x080F
        "00101010", -- 0x0810
        "00000010", -- 0x0811
        "00001000", -- 0x0812
        "10010101", -- 0x0813
        "00010010", -- 0x0814
        "00100000", -- 0x0815
        "10110011", -- 0x0816
        "00010010", -- 0x0817
        "00010100", -- 0x0818
        "11011100", -- 0x0819
        "01110100", -- 0x081A
        "01111001", -- 0x081B
        "00010010", -- 0x081C
        "00100000", -- 0x081D
        "01110111", -- 0x081E
        "10000000", -- 0x081F
        "01110100", -- 0x0820
        "00010010", -- 0x0821
        "00100010", -- 0x0822
        "01111100", -- 0x0823
        "01110100", -- 0x0824
        "00001011", -- 0x0825
        "11110000", -- 0x0826
        "10100011", -- 0x0827
        "01110100", -- 0x0828
        "10001001", -- 0x0829
        "11110000", -- 0x082A
        "10100011", -- 0x082B
        "11100100", -- 0x082C
        "00010010", -- 0x082D
        "00100010", -- 0x082E
        "10111110", -- 0x082F
        "01110100", -- 0x0830
        "01100110", -- 0x0831
        "11110000", -- 0x0832
        "10100011", -- 0x0833
        "00010010", -- 0x0834
        "00100011", -- 0x0835
        "10001111", -- 0x0836
        "00010010", -- 0x0837
        "00010100", -- 0x0838
        "11011100", -- 0x0839
        "01110100", -- 0x083A
        "01111010", -- 0x083B
        "00010010", -- 0x083C
        "00100000", -- 0x083D
        "01110111", -- 0x083E
        "10000000", -- 0x083F
        "01010100", -- 0x0840
        "00010010", -- 0x0841
        "00100011", -- 0x0842
        "00011110", -- 0x0843
        "01110100", -- 0x0844
        "00001110", -- 0x0845
        "11110000", -- 0x0846
        "10100011", -- 0x0847
        "01110100", -- 0x0848
        "00000001", -- 0x0849
        "11110000", -- 0x084A
        "10010000", -- 0x084B
        "00011000", -- 0x084C
        "00001010", -- 0x084D
        "01110100", -- 0x084E
        "11110100", -- 0x084F
        "00010010", -- 0x0850
        "00100011", -- 0x0851
        "10000001", -- 0x0852
        "01110100", -- 0x0853
        "00001001", -- 0x0854
        "11110000", -- 0x0855
        "00010010", -- 0x0856
        "00100011", -- 0x0857
        "11001110", -- 0x0858
        "01110100", -- 0x0859
        "00110010", -- 0x085A
        "00010010", -- 0x085B
        "00100011", -- 0x085C
        "10000001", -- 0x085D
        "01110100", -- 0x085E
        "00001111", -- 0x085F
        "11110000", -- 0x0860
        "00010010", -- 0x0861
        "00100011", -- 0x0862
        "11001110", -- 0x0863
        "11100100", -- 0x0864
        "00010010", -- 0x0865
        "00100011", -- 0x0866
        "10000001", -- 0x0867
        "00010010", -- 0x0868
        "00100100", -- 0x0869
        "01111101", -- 0x086A
        "01111000", -- 0x086B
        "00000000", -- 0x086C
        "10000000", -- 0x086D
        "00100110", -- 0x086E
        "00010010", -- 0x086F
        "00100010", -- 0x0870
        "01111100", -- 0x0871
        "01110100", -- 0x0872
        "10100000", -- 0x0873
        "11110000", -- 0x0874
        "10100011", -- 0x0875
        "01110100", -- 0x0876
        "00000010", -- 0x0877
        "11110000", -- 0x0878
        "10100011", -- 0x0879
        "01110100", -- 0x087A
        "01011000", -- 0x087B
        "00010010", -- 0x087C
        "00100011", -- 0x087D
        "10010110", -- 0x087E
        "11100100", -- 0x087F
        "11110000", -- 0x0880
        "10100011", -- 0x0881
        "01110100", -- 0x0882
        "01100100", -- 0x0883
        "00010010", -- 0x0884
        "00100001", -- 0x0885
        "11010100", -- 0x0886
        "01110100", -- 0x0887
        "00001010", -- 0x0888
        "00010010", -- 0x0889
        "00100011", -- 0x088A
        "00010110", -- 0x088B
        "11100100", -- 0x088C
        "11110000", -- 0x088D
        "00010010", -- 0x088E
        "00100100", -- 0x088F
        "00101010", -- 0x0890
        "10000000", -- 0x0891
        "00000010", -- 0x0892
        "01111000", -- 0x0893
        "11001100", -- 0x0894
        "11101000", -- 0x0895
        "00100010", -- 0x0896
        "10010000", -- 0x0897
        "00000000", -- 0x0898
        "00000011", -- 0x0899
        "11100000", -- 0x089A
        "10110100", -- 0x089B
        "00010101", -- 0x089C
        "00001101", -- 0x089D
        "10010000", -- 0x089E
        "00000000", -- 0x089F
        "00000000", -- 0x08A0
        "11100000", -- 0x08A1
        "10010000", -- 0x08A2
        "00000000", -- 0x08A3
        "00000010", -- 0x08A4
        "11110000", -- 0x08A5
        "10010000", -- 0x08A6
        "00000000", -- 0x08A7
        "00000011", -- 0x08A8
        "11100100", -- 0x08A9
        "11110000", -- 0x08AA
        "10010000", -- 0x08AB
        "00000000", -- 0x08AC
        "00000100", -- 0x08AD
        "11100000", -- 0x08AE
        "01100000", -- 0x08AF
        "00000011", -- 0x08B0
        "00000010", -- 0x08B1
        "00001001", -- 0x08B2
        "10000000", -- 0x08B3
        "10010000", -- 0x08B4
        "00000000", -- 0x08B5
        "00000100", -- 0x08B6
        "01110100", -- 0x08B7
        "00000001", -- 0x08B8
        "11110000", -- 0x08B9
        "00010010", -- 0x08BA
        "00100000", -- 0x08BB
        "11001111", -- 0x08BC
        "01000000", -- 0x08BD
        "00000101", -- 0x08BE
        "00010010", -- 0x08BF
        "00100000", -- 0x08C0
        "11001111", -- 0x08C1
        "10000000", -- 0x08C2
        "00010001", -- 0x08C3
        "10010000", -- 0x08C4
        "00000000", -- 0x08C5
        "00000010", -- 0x08C6
        "11100000", -- 0x08C7
        "11111000", -- 0x08C8
        "01111011", -- 0x08C9
        "00100100", -- 0x08CA
        "11101011", -- 0x08CB
        "11000011", -- 0x08CC
        "10011000", -- 0x08CD
        "11111001", -- 0x08CE
        "10010000", -- 0x08CF
        "00000000", -- 0x08D0
        "00000000", -- 0x08D1
        "11100000", -- 0x08D2
        "11111010", -- 0x08D3
        "00101001", -- 0x08D4
        "11111001", -- 0x08D5
        "10010000", -- 0x08D6
        "00000001", -- 0x08D7
        "00011000", -- 0x08D8
        "11101001", -- 0x08D9
        "11110000", -- 0x08DA
        "11101001", -- 0x08DB
        "11111000", -- 0x08DC
        "11010011", -- 0x08DD
        "10010100", -- 0x08DE
        "00000010", -- 0x08DF
        "01010000", -- 0x08E0
        "00000011", -- 0x08E1
        "00000010", -- 0x08E2
        "00001001", -- 0x08E3
        "01111011", -- 0x08E4
        "00010010", -- 0x08E5
        "00100000", -- 0x08E6
        "00101001", -- 0x08E7
        "11100000", -- 0x08E8
        "10110100", -- 0x08E9
        "00011110", -- 0x08EA
        "01010101", -- 0x08EB
        "11101000", -- 0x08EC
        "11010011", -- 0x08ED
        "10010100", -- 0x08EE
        "00000100", -- 0x08EF
        "01010000", -- 0x08F0
        "00000011", -- 0x08F1
        "00000010", -- 0x08F2
        "00001001", -- 0x08F3
        "01111011", -- 0x08F4
        "00010010", -- 0x08F5
        "00011101", -- 0x08F6
        "01010001", -- 0x08F7
        "00010010", -- 0x08F8
        "00100100", -- 0x08F9
        "00011110", -- 0x08FA
        "11111111", -- 0x08FB
        "11100100", -- 0x08FC
        "00111000", -- 0x08FD
        "11111110", -- 0x08FE
        "00010010", -- 0x08FF
        "00100000", -- 0x0900
        "10000110", -- 0x0901
        "10010000", -- 0x0902
        "00011000", -- 0x0903
        "00100011", -- 0x0904
        "11110000", -- 0x0905
        "00010010", -- 0x0906
        "00100011", -- 0x0907
        "10110010", -- 0x0908
        "00100100", -- 0x0909
        "00000100", -- 0x090A
        "11111111", -- 0x090B
        "11100100", -- 0x090C
        "00111000", -- 0x090D
        "11111110", -- 0x090E
        "00010010", -- 0x090F
        "00100000", -- 0x0910
        "10000110", -- 0x0911
        "10010000", -- 0x0912
        "00011000", -- 0x0913
        "00100100", -- 0x0914
        "11110000", -- 0x0915
        "11100000", -- 0x0916
        "11110101", -- 0x0917
        "00010100", -- 0x0918
        "01111100", -- 0x0919
        "00000000", -- 0x091A
        "01111101", -- 0x091B
        "00000100", -- 0x091C
        "01111110", -- 0x091D
        "00011000", -- 0x091E
        "01111111", -- 0x091F
        "00100000", -- 0x0920
        "00010010", -- 0x0921
        "00010111", -- 0x0922
        "10001110", -- 0x0923
        "10110101", -- 0x0924
        "00010100", -- 0x0925
        "00000010", -- 0x0926
        "10000000", -- 0x0927
        "00000011", -- 0x0928
        "00000010", -- 0x0929
        "00001001", -- 0x092A
        "00110101", -- 0x092B
        "01111110", -- 0x092C
        "00011000", -- 0x092D
        "01111111", -- 0x092E
        "00100000", -- 0x092F
        "00010010", -- 0x0930
        "00010010", -- 0x0931
        "01100111", -- 0x0932
        "10000000", -- 0x0933
        "00000101", -- 0x0934
        "01111111", -- 0x0935
        "00010101", -- 0x0936
        "00010010", -- 0x0937
        "00011000", -- 0x0938
        "01010010", -- 0x0939
        "00010010", -- 0x093A
        "00100011", -- 0x093B
        "10110010", -- 0x093C
        "00100100", -- 0x093D
        "00000101", -- 0x093E
        "10000000", -- 0x093F
        "00101101", -- 0x0940
        "00010010", -- 0x0941
        "00100000", -- 0x0942
        "00101001", -- 0x0943
        "00010010", -- 0x0944
        "00011101", -- 0x0945
        "01010001", -- 0x0946
        "11100000", -- 0x0947
        "11110101", -- 0x0948
        "00010100", -- 0x0949
        "01111100", -- 0x094A
        "00000000", -- 0x094B
        "01111101", -- 0x094C
        "00000010", -- 0x094D
        "01111110", -- 0x094E
        "00011000", -- 0x094F
        "01111111", -- 0x0950
        "00100000", -- 0x0951
        "00010010", -- 0x0952
        "00010111", -- 0x0953
        "10001110", -- 0x0954
        "10110101", -- 0x0955
        "00010100", -- 0x0956
        "00000010", -- 0x0957
        "10000000", -- 0x0958
        "00000011", -- 0x0959
        "00000010", -- 0x095A
        "00001001", -- 0x095B
        "01100110", -- 0x095C
        "01111110", -- 0x095D
        "00011000", -- 0x095E
        "01111111", -- 0x095F
        "00100000", -- 0x0960
        "00010010", -- 0x0961
        "00001101", -- 0x0962
        "01010011", -- 0x0963
        "10000000", -- 0x0964
        "00000101", -- 0x0965
        "01111111", -- 0x0966
        "00010101", -- 0x0967
        "00010010", -- 0x0968
        "00011000", -- 0x0969
        "01010010", -- 0x096A
        "00010010", -- 0x096B
        "00100100", -- 0x096C
        "00011110", -- 0x096D
        "11111111", -- 0x096E
        "11101000", -- 0x096F
        "00110100", -- 0x0970
        "00000000", -- 0x0971
        "11111110", -- 0x0972
        "00010010", -- 0x0973
        "00100011", -- 0x0974
        "11110001", -- 0x0975
        "10010000", -- 0x0976
        "00000000", -- 0x0977
        "00000010", -- 0x0978
        "11101101", -- 0x0979
        "11110000", -- 0x097A
        "10010000", -- 0x097B
        "00000000", -- 0x097C
        "00000100", -- 0x097D
        "11100100", -- 0x097E
        "11110000", -- 0x097F
        "00100010", -- 0x0980
        "00010010", -- 0x0981
        "00011100", -- 0x0982
        "01100100", -- 0x0983
        "10000000", -- 0x0984
        "01010000", -- 0x0985
        "11100000", -- 0x0986
        "11000000", -- 0x0987
        "11100000", -- 0x0988
        "10100011", -- 0x0989
        "11100000", -- 0x098A
        "11000000", -- 0x098B
        "11100000", -- 0x098C
        "10100011", -- 0x098D
        "11100000", -- 0x098E
        "11000000", -- 0x098F
        "11100000", -- 0x0990
        "10100011", -- 0x0991
        "11100000", -- 0x0992
        "11000000", -- 0x0993
        "11100000", -- 0x0994
        "10000000", -- 0x0995
        "00111111", -- 0x0996
        "11100100", -- 0x0997
        "10010011", -- 0x0998
        "11000000", -- 0x0999
        "11100000", -- 0x099A
        "10100011", -- 0x099B
        "11100100", -- 0x099C
        "10010011", -- 0x099D
        "11000000", -- 0x099E
        "11100000", -- 0x099F
        "10100011", -- 0x09A0
        "11100100", -- 0x09A1
        "10010011", -- 0x09A2
        "11000000", -- 0x09A3
        "11100000", -- 0x09A4
        "10100011", -- 0x09A5
        "11100100", -- 0x09A6
        "10010011", -- 0x09A7
        "11000000", -- 0x09A8
        "11100000", -- 0x09A9
        "10000000", -- 0x09AA
        "00101010", -- 0x09AB
        "10001000", -- 0x09AC
        "11110000", -- 0x09AD
        "11100110", -- 0x09AE
        "11000000", -- 0x09AF
        "11100000", -- 0x09B0
        "00001000", -- 0x09B1
        "11100110", -- 0x09B2
        "11000000", -- 0x09B3
        "11100000", -- 0x09B4
        "00001000", -- 0x09B5
        "11100110", -- 0x09B6
        "11000000", -- 0x09B7
        "11100000", -- 0x09B8
        "00001000", -- 0x09B9
        "11100110", -- 0x09BA
        "11000000", -- 0x09BB
        "11100000", -- 0x09BC
        "10101000", -- 0x09BD
        "11110000", -- 0x09BE
        "10000000", -- 0x09BF
        "00010101", -- 0x09C0
        "10001000", -- 0x09C1
        "11110000", -- 0x09C2
        "11100010", -- 0x09C3
        "11000000", -- 0x09C4
        "11100000", -- 0x09C5
        "00001000", -- 0x09C6
        "11100010", -- 0x09C7
        "11000000", -- 0x09C8
        "11100000", -- 0x09C9
        "00001000", -- 0x09CA
        "11100010", -- 0x09CB
        "11000000", -- 0x09CC
        "11100000", -- 0x09CD
        "00001000", -- 0x09CE
        "11100010", -- 0x09CF
        "11000000", -- 0x09D0
        "11100000", -- 0x09D1
        "10101000", -- 0x09D2
        "11110000", -- 0x09D3
        "10000000", -- 0x09D4
        "00000000", -- 0x09D5
        "11100100", -- 0x09D6
        "11000000", -- 0x09D7
        "11100000", -- 0x09D8
        "11000000", -- 0x09D9
        "11100000", -- 0x09DA
        "11000000", -- 0x09DB
        "11100000", -- 0x09DC
        "11000000", -- 0x09DD
        "11100000", -- 0x09DE
        "11100101", -- 0x09DF
        "10000001", -- 0x09E0
        "11001011", -- 0x09E1
        "11000000", -- 0x09E2
        "11100000", -- 0x09E3
        "11101010", -- 0x09E4
        "11000000", -- 0x09E5
        "11100000", -- 0x09E6
        "11101001", -- 0x09E7
        "11000000", -- 0x09E8
        "11100000", -- 0x09E9
        "01110100", -- 0x09EA
        "11111100", -- 0x09EB
        "00101011", -- 0x09EC
        "11001000", -- 0x09ED
        "11000000", -- 0x09EE
        "11100000", -- 0x09EF
        "01111010", -- 0x09F0
        "00000100", -- 0x09F1
        "11101111", -- 0x09F2
        "00010010", -- 0x09F3
        "00001010", -- 0x09F4
        "01001111", -- 0x09F5
        "00011011", -- 0x09F6
        "11101110", -- 0x09F7
        "00010010", -- 0x09F8
        "00001010", -- 0x09F9
        "01000101", -- 0x09FA
        "00011011", -- 0x09FB
        "11101101", -- 0x09FC
        "00010010", -- 0x09FD
        "00001010", -- 0x09FE
        "01001001", -- 0x09FF
        "00011011", -- 0x0A00
        "11101100", -- 0x0A01
        "00010010", -- 0x0A02
        "00001010", -- 0x0A03
        "01001101", -- 0x0A04
        "00011000", -- 0x0A05
        "00001011", -- 0x0A06
        "00001011", -- 0x0A07
        "11101111", -- 0x0A08
        "00010010", -- 0x0A09
        "00001010", -- 0x0A0A
        "01000101", -- 0x0A0B
        "00011011", -- 0x0A0C
        "11101110", -- 0x0A0D
        "00010010", -- 0x0A0E
        "00001010", -- 0x0A0F
        "01001001", -- 0x0A10
        "00011011", -- 0x0A11
        "11101101", -- 0x0A12
        "00010010", -- 0x0A13
        "00001010", -- 0x0A14
        "01001101", -- 0x0A15
        "00011000", -- 0x0A16
        "00001011", -- 0x0A17
        "11101111", -- 0x0A18
        "00010010", -- 0x0A19
        "00001010", -- 0x0A1A
        "01001001", -- 0x0A1B
        "00011011", -- 0x0A1C
        "11101110", -- 0x0A1D
        "00010010", -- 0x0A1E
        "00001010", -- 0x0A1F
        "01001101", -- 0x0A20
        "00011000", -- 0x0A21
        "11101111", -- 0x0A22
        "00010010", -- 0x0A23
        "00001010", -- 0x0A24
        "01001101", -- 0x0A25
        "11010000", -- 0x0A26
        "11100000", -- 0x0A27
        "11111000", -- 0x0A28
        "11010000", -- 0x0A29
        "11100000", -- 0x0A2A
        "11111001", -- 0x0A2B
        "11010000", -- 0x0A2C
        "11100000", -- 0x0A2D
        "11111010", -- 0x0A2E
        "11010000", -- 0x0A2F
        "11100000", -- 0x0A30
        "11111011", -- 0x0A31
        "11010000", -- 0x0A32
        "11100000", -- 0x0A33
        "11111111", -- 0x0A34
        "11010000", -- 0x0A35
        "11100000", -- 0x0A36
        "11111110", -- 0x0A37
        "11010000", -- 0x0A38
        "11100000", -- 0x0A39
        "11111101", -- 0x0A3A
        "11010000", -- 0x0A3B
        "11100000", -- 0x0A3C
        "11111100", -- 0x0A3D
        "11100101", -- 0x0A3E
        "10000001", -- 0x0A3F
        "00100100", -- 0x0A40
        "11111100", -- 0x0A41
        "11110101", -- 0x0A42
        "10000001", -- 0x0A43
        "00100010", -- 0x0A44
        "01111010", -- 0x0A45
        "00000011", -- 0x0A46
        "10000000", -- 0x0A47
        "00000110", -- 0x0A48
        "01111010", -- 0x0A49
        "00000010", -- 0x0A4A
        "10000000", -- 0x0A4B
        "00000010", -- 0x0A4C
        "01111010", -- 0x0A4D
        "00000001", -- 0x0A4E
        "11110101", -- 0x0A4F
        "11110000", -- 0x0A50
        "11101011", -- 0x0A51
        "11111001", -- 0x0A52
        "11100110", -- 0x0A53
        "10100100", -- 0x0A54
        "00100111", -- 0x0A55
        "11110111", -- 0x0A56
        "11011010", -- 0x0A57
        "00000001", -- 0x0A58
        "00100010", -- 0x0A59
        "11100101", -- 0x0A5A
        "11110000", -- 0x0A5B
        "00011001", -- 0x0A5C
        "00110111", -- 0x0A5D
        "11110111", -- 0x0A5E
        "11011010", -- 0x0A5F
        "00000001", -- 0x0A60
        "00100010", -- 0x0A61
        "01010000", -- 0x0A62
        "00000110", -- 0x0A63
        "00011001", -- 0x0A64
        "11100100", -- 0x0A65
        "00110111", -- 0x0A66
        "11110111", -- 0x0A67
        "11011010", -- 0x0A68
        "11111000", -- 0x0A69
        "00100010", -- 0x0A6A
        "10010000", -- 0x0A6B
        "00000001", -- 0x0A6C
        "10001101", -- 0x0A6D
        "11100101", -- 0x0A6E
        "11001101", -- 0x0A6F
        "11110000", -- 0x0A70
        "10100011", -- 0x0A71
        "11100101", -- 0x0A72
        "11000101", -- 0x0A73
        "11110000", -- 0x0A74
        "10010000", -- 0x0A75
        "00000001", -- 0x0A76
        "10010000", -- 0x0A77
        "11100101", -- 0x0A78
        "10111101", -- 0x0A79
        "11110000", -- 0x0A7A
        "10010000", -- 0x0A7B
        "00000001", -- 0x0A7C
        "10001111", -- 0x0A7D
        "11100101", -- 0x0A7E
        "10010101", -- 0x0A7F
        "11110000", -- 0x0A80
        "10100011", -- 0x0A81
        "10100011", -- 0x0A82
        "11100101", -- 0x0A83
        "10100101", -- 0x0A84
        "11110000", -- 0x0A85
        "10010000", -- 0x0A86
        "00000001", -- 0x0A87
        "10010010", -- 0x0A88
        "11100101", -- 0x0A89
        "10011101", -- 0x0A8A
        "11110000", -- 0x0A8B
        "11100101", -- 0x0A8C
        "10011101", -- 0x0A8D
        "11111101", -- 0x0A8E
        "11100100", -- 0x0A8F
        "11111110", -- 0x0A90
        "01111100", -- 0x0A91
        "00000000", -- 0x0A92
        "01111111", -- 0x0A93
        "11111111", -- 0x0A94
        "00010010", -- 0x0A95
        "00011110", -- 0x0A96
        "10110110", -- 0x0A97
        "11100101", -- 0x0A98
        "10100101", -- 0x0A99
        "11000011", -- 0x0A9A
        "00010011", -- 0x0A9B
        "11111000", -- 0x0A9C
        "00101111", -- 0x0A9D
        "11111111", -- 0x0A9E
        "11100100", -- 0x0A9F
        "00111110", -- 0x0AA0
        "11111110", -- 0x0AA1
        "11100101", -- 0x0AA2
        "10100101", -- 0x0AA3
        "11111101", -- 0x0AA4
        "01111100", -- 0x0AA5
        "00000000", -- 0x0AA6
        "00010010", -- 0x0AA7
        "00001111", -- 0x0AA8
        "11010100", -- 0x0AA9
        "11101111", -- 0x0AAA
        "10010000", -- 0x0AAB
        "00000000", -- 0x0AAC
        "00011000", -- 0x0AAD
        "00010010", -- 0x0AAE
        "00100010", -- 0x0AAF
        "11101011", -- 0x0AB0
        "11100000", -- 0x0AB1
        "10010000", -- 0x0AB2
        "00000001", -- 0x0AB3
        "10010110", -- 0x0AB4
        "11110000", -- 0x0AB5
        "11100000", -- 0x0AB6
        "00100100", -- 0x0AB7
        "00101001", -- 0x0AB8
        "10100011", -- 0x0AB9
        "11110000", -- 0x0ABA
        "00010010", -- 0x0ABB
        "00100000", -- 0x0ABC
        "11011101", -- 0x0ABD
        "11100100", -- 0x0ABE
        "11111010", -- 0x0ABF
        "11100100", -- 0x0AC0
        "11111011", -- 0x0AC1
        "00100000", -- 0x0AC2
        "10100001", -- 0x0AC3
        "00000110", -- 0x0AC4
        "11100101", -- 0x0AC5
        "10100000", -- 0x0AC6
        "01010100", -- 0x0AC7
        "00000101", -- 0x0AC8
        "01100000", -- 0x0AC9
        "00000110", -- 0x0ACA
        "00100000", -- 0x0ACB
        "10100001", -- 0x0ACC
        "00000101", -- 0x0ACD
        "00100000", -- 0x0ACE
        "10100101", -- 0x0ACF
        "00000010", -- 0x0AD0
        "01111011", -- 0x0AD1
        "00000001", -- 0x0AD2
        "11101011", -- 0x0AD3
        "01110000", -- 0x0AD4
        "00000110", -- 0x0AD5
        "00100000", -- 0x0AD6
        "10100001", -- 0x0AD7
        "00000101", -- 0x0AD8
        "00100000", -- 0x0AD9
        "10100101", -- 0x0ADA
        "00000010", -- 0x0ADB
        "01111010", -- 0x0ADC
        "00000001", -- 0x0ADD
        "11100100", -- 0x0ADE
        "11111011", -- 0x0ADF
        "11100100", -- 0x0AE0
        "11111100", -- 0x0AE1
        "00100000", -- 0x0AE2
        "10100000", -- 0x0AE3
        "00000101", -- 0x0AE4
        "00100000", -- 0x0AE5
        "10100010", -- 0x0AE6
        "00000010", -- 0x0AE7
        "01111100", -- 0x0AE8
        "00000001", -- 0x0AE9
        "11101100", -- 0x0AEA
        "01110000", -- 0x0AEB
        "00001100", -- 0x0AEC
        "00100000", -- 0x0AED
        "10100000", -- 0x0AEE
        "00000011", -- 0x0AEF
        "00110000", -- 0x0AF0
        "10100100", -- 0x0AF1
        "00000110", -- 0x0AF2
        "00100000", -- 0x0AF3
        "10100010", -- 0x0AF4
        "00000101", -- 0x0AF5
        "00100000", -- 0x0AF6
        "10100100", -- 0x0AF7
        "00000010", -- 0x0AF8
        "01111011", -- 0x0AF9
        "00000001", -- 0x0AFA
        "11100101", -- 0x0AFB
        "11101101", -- 0x0AFC
        "00010010", -- 0x0AFD
        "00100010", -- 0x0AFE
        "01101000", -- 0x0AFF
        "11111100", -- 0x0B00
        "11101011", -- 0x0B01
        "00100101", -- 0x0B02
        "11100000", -- 0x0B03
        "11111011", -- 0x0B04
        "11101010", -- 0x0B05
        "00100011", -- 0x0B06
        "00100011", -- 0x0B07
        "01010100", -- 0x0B08
        "11111100", -- 0x0B09
        "11111010", -- 0x0B0A
        "11100101", -- 0x0B0B
        "11101101", -- 0x0B0C
        "00010010", -- 0x0B0D
        "00100010", -- 0x0B0E
        "01011110", -- 0x0B0F
        "11000100", -- 0x0B10
        "00000011", -- 0x0B11
        "01010100", -- 0x0B12
        "11111000", -- 0x0B13
        "11111101", -- 0x0B14
        "10010000", -- 0x0B15
        "00000001", -- 0x0B16
        "00011011", -- 0x0B17
        "11100000", -- 0x0B18
        "11000100", -- 0x0B19
        "00100011", -- 0x0B1A
        "01010100", -- 0x0B1B
        "11100000", -- 0x0B1C
        "11111110", -- 0x0B1D
        "11101001", -- 0x0B1E
        "00000011", -- 0x0B1F
        "00000011", -- 0x0B20
        "01010100", -- 0x0B21
        "11000000", -- 0x0B22
        "11111001", -- 0x0B23
        "11101000", -- 0x0B24
        "00000011", -- 0x0B25
        "01010100", -- 0x0B26
        "10000000", -- 0x0B27
        "01001001", -- 0x0B28
        "01001110", -- 0x0B29
        "01001101", -- 0x0B2A
        "01001010", -- 0x0B2B
        "01001011", -- 0x0B2C
        "01001100", -- 0x0B2D
        "10010000", -- 0x0B2E
        "00000001", -- 0x0B2F
        "10011000", -- 0x0B30
        "11110000", -- 0x0B31
        "00100010", -- 0x0B32
        "11101111", -- 0x0B33
        "01100000", -- 0x0B34
        "00010001", -- 0x0B35
        "00010100", -- 0x0B36
        "01100000", -- 0x0B37
        "01001000", -- 0x0B38
        "00100100", -- 0x0B39
        "11111110", -- 0x0B3A
        "01100000", -- 0x0B3B
        "01111101", -- 0x0B3C
        "00100100", -- 0x0B3D
        "11111100", -- 0x0B3E
        "01110000", -- 0x0B3F
        "00000011", -- 0x0B40
        "00000010", -- 0x0B41
        "00001011", -- 0x0B42
        "11010110", -- 0x0B43
        "00000010", -- 0x0B44
        "00001011", -- 0x0B45
        "11100110", -- 0x0B46
        "00010010", -- 0x0B47
        "00100010", -- 0x0B48
        "10011010", -- 0x0B49
        "10010000", -- 0x0B4A
        "00000001", -- 0x0B4B
        "00011011", -- 0x0B4C
        "11100100", -- 0x0B4D
        "11110000", -- 0x0B4E
        "10010000", -- 0x0B4F
        "00000000", -- 0x0B50
        "00010000", -- 0x0B51
        "11100100", -- 0x0B52
        "11110000", -- 0x0B53
        "10100011", -- 0x0B54
        "01110100", -- 0x0B55
        "11111111", -- 0x0B56
        "11110000", -- 0x0B57
        "11100100", -- 0x0B58
        "11111101", -- 0x0B59
        "11111100", -- 0x0B5A
        "00010010", -- 0x0B5B
        "00100011", -- 0x0B5C
        "01011110", -- 0x0B5D
        "00010010", -- 0x0B5E
        "00100100", -- 0x0B5F
        "01001110", -- 0x0B60
        "11100100", -- 0x0B61
        "11111101", -- 0x0B62
        "11111100", -- 0x0B63
        "01111110", -- 0x0B64
        "00011010", -- 0x0B65
        "01111111", -- 0x0B66
        "00101011", -- 0x0B67
        "00010010", -- 0x0B68
        "00010100", -- 0x0B69
        "00010100", -- 0x0B6A
        "01111100", -- 0x0B6B
        "00001111", -- 0x0B6C
        "01111101", -- 0x0B6D
        "10100000", -- 0x0B6E
        "01111110", -- 0x0B6F
        "00001111", -- 0x0B70
        "01111111", -- 0x0B71
        "00111001", -- 0x0B72
        "00010010", -- 0x0B73
        "00010100", -- 0x0B74
        "00010100", -- 0x0B75
        "00010010", -- 0x0B76
        "00100010", -- 0x0B77
        "10100011", -- 0x0B78
        "00010010", -- 0x0B79
        "00100010", -- 0x0B7A
        "10101100", -- 0x0B7B
        "00010010", -- 0x0B7C
        "00100100", -- 0x0B7D
        "10011101", -- 0x0B7E
        "10000000", -- 0x0B7F
        "01101000", -- 0x0B80
        "00010010", -- 0x0B81
        "00100010", -- 0x0B82
        "10011010", -- 0x0B83
        "10010000", -- 0x0B84
        "00000001", -- 0x0B85
        "00011100", -- 0x0B86
        "01110100", -- 0x0B87
        "00000001", -- 0x0B88
        "11110000", -- 0x0B89
        "10010000", -- 0x0B8A
        "00000001", -- 0x0B8B
        "10010011", -- 0x0B8C
        "00010010", -- 0x0B8D
        "00100011", -- 0x0B8E
        "01000110", -- 0x0B8F
        "10010000", -- 0x0B90
        "00000001", -- 0x0B91
        "01000110", -- 0x0B92
        "00010010", -- 0x0B93
        "00011011", -- 0x0B94
        "11010001", -- 0x0B95
        "00010010", -- 0x0B96
        "00011001", -- 0x0B97
        "01001000", -- 0x0B98
        "10010000", -- 0x0B99
        "00000001", -- 0x0B9A
        "01001010", -- 0x0B9B
        "00010010", -- 0x0B9C
        "00011011", -- 0x0B9D
        "11010001", -- 0x0B9E
        "01111100", -- 0x0B9F
        "00000000", -- 0x0BA0
        "01111101", -- 0x0BA1
        "00001010", -- 0x0BA2
        "01111110", -- 0x0BA3
        "00000001", -- 0x0BA4
        "01111111", -- 0x0BA5
        "01000110", -- 0x0BA6
        "00010010", -- 0x0BA7
        "00010111", -- 0x0BA8
        "10001110", -- 0x0BA9
        "10010000", -- 0x0BAA
        "00000001", -- 0x0BAB
        "01010000", -- 0x0BAC
        "11110000", -- 0x0BAD
        "00010010", -- 0x0BAE
        "00100100", -- 0x0BAF
        "10011101", -- 0x0BB0
        "01111101", -- 0x0BB1
        "00001011", -- 0x0BB2
        "01111110", -- 0x0BB3
        "00000001", -- 0x0BB4
        "01111111", -- 0x0BB5
        "01000110", -- 0x0BB6
        "00000010", -- 0x0BB7
        "00011011", -- 0x0BB8
        "10101011", -- 0x0BB9
        "00010010", -- 0x0BBA
        "00100011", -- 0x0BBB
        "11100011", -- 0x0BBC
        "01110101", -- 0x0BBD
        "11100101", -- 0x0BBE
        "11111111", -- 0x0BBF
        "11100100", -- 0x0BC0
        "11111110", -- 0x0BC1
        "11111101", -- 0x0BC2
        "11111100", -- 0x0BC3
        "01111111", -- 0x0BC4
        "01100100", -- 0x0BC5
        "00010010", -- 0x0BC6
        "00010110", -- 0x0BC7
        "00110100", -- 0x0BC8
        "01110101", -- 0x0BC9
        "11100101", -- 0x0BCA
        "01111010", -- 0x0BCB
        "01110101", -- 0x0BCC
        "10110000", -- 0x0BCD
        "00000000", -- 0x0BCE
        "10010000", -- 0x0BCF
        "00000001", -- 0x0BD0
        "00011100", -- 0x0BD1
        "01110100", -- 0x0BD2
        "00000011", -- 0x0BD3
        "10000000", -- 0x0BD4
        "00010111", -- 0x0BD5
        "00010010", -- 0x0BD6
        "00100011", -- 0x0BD7
        "11100011", -- 0x0BD8
        "00010010", -- 0x0BD9
        "00100010", -- 0x0BDA
        "01010100", -- 0x0BDB
        "00010010", -- 0x0BDC
        "00011111", -- 0x0BDD
        "01101100", -- 0x0BDE
        "10010000", -- 0x0BDF
        "00000001", -- 0x0BE0
        "00011100", -- 0x0BE1
        "01110100", -- 0x0BE2
        "00000111", -- 0x0BE3
        "10000000", -- 0x0BE4
        "00000111", -- 0x0BE5
        "00010010", -- 0x0BE6
        "00100010", -- 0x0BE7
        "10011010", -- 0x0BE8
        "10010000", -- 0x0BE9
        "00000001", -- 0x0BEA
        "00011100", -- 0x0BEB
        "11100100", -- 0x0BEC
        "11110000", -- 0x0BED
        "00100010", -- 0x0BEE
        "01110101", -- 0x0BEF
        "10100000", -- 0x0BF0
        "00000001", -- 0x0BF1
        "00010010", -- 0x0BF2
        "00011110", -- 0x0BF3
        "11100000", -- 0x0BF4
        "01111100", -- 0x0BF5
        "00000000", -- 0x0BF6
        "01111101", -- 0x0BF7
        "01100100", -- 0x0BF8
        "01111110", -- 0x0BF9
        "00001000", -- 0x0BFA
        "01111111", -- 0x0BFB
        "10010111", -- 0x0BFC
        "00010010", -- 0x0BFD
        "00100011", -- 0x0BFE
        "10111001", -- 0x0BFF
        "01111110", -- 0x0C00
        "00001111", -- 0x0C01
        "01111111", -- 0x0C02
        "00111001", -- 0x0C03
        "00010010", -- 0x0C04
        "00010001", -- 0x0C05
        "00000010", -- 0x0C06
        "01111100", -- 0x0C07
        "00000001", -- 0x0C08
        "01111101", -- 0x0C09
        "11110100", -- 0x0C0A
        "01111110", -- 0x0C0B
        "00001010", -- 0x0C0C
        "01111111", -- 0x0C0D
        "01101011", -- 0x0C0E
        "00010010", -- 0x0C0F
        "00100011", -- 0x0C10
        "10111001", -- 0x0C11
        "01111110", -- 0x0C12
        "00000011", -- 0x0C13
        "01111111", -- 0x0C14
        "00101010", -- 0x0C15
        "00010010", -- 0x0C16
        "00100011", -- 0x0C17
        "10111001", -- 0x0C18
        "01111110", -- 0x0C19
        "00011010", -- 0x0C1A
        "01111111", -- 0x0C1B
        "00101011", -- 0x0C1C
        "00010010", -- 0x0C1D
        "00100011", -- 0x0C1E
        "10111001", -- 0x0C1F
        "01111110", -- 0x0C20
        "00000100", -- 0x0C21
        "01111111", -- 0x0C22
        "11001101", -- 0x0C23
        "00010010", -- 0x0C24
        "00010001", -- 0x0C25
        "00000010", -- 0x0C26
        "01111111", -- 0x0C27
        "00000000", -- 0x0C28
        "00010010", -- 0x0C29
        "00001011", -- 0x0C2A
        "00110011", -- 0x0C2B
        "00010010", -- 0x0C2C
        "00100001", -- 0x0C2D
        "00111000", -- 0x0C2E
        "00010010", -- 0x0C2F
        "00010011", -- 0x0C30
        "10101101", -- 0x0C31
        "01110101", -- 0x0C32
        "10100000", -- 0x0C33
        "00000001", -- 0x0C34
        "01110101", -- 0x0C35
        "10100000", -- 0x0C36
        "00000010", -- 0x0C37
        "11100101", -- 0x0C38
        "10011011", -- 0x0C39
        "01010100", -- 0x0C3A
        "00000001", -- 0x0C3B
        "01100000", -- 0x0C3C
        "00101110", -- 0x0C3D
        "11100101", -- 0x0C3E
        "10001011", -- 0x0C3F
        "11111001", -- 0x0C40
        "01111000", -- 0x0C41
        "00000000", -- 0x0C42
        "10010000", -- 0x0C43
        "00000001", -- 0x0C44
        "00100011", -- 0x0C45
        "11101000", -- 0x0C46
        "11110000", -- 0x0C47
        "11101001", -- 0x0C48
        "10100011", -- 0x0C49
        "11110000", -- 0x0C4A
        "10010000", -- 0x0C4B
        "00000001", -- 0x0C4C
        "00100011", -- 0x0C4D
        "01111111", -- 0x0C4E
        "00001000", -- 0x0C4F
        "00010010", -- 0x0C50
        "00011110", -- 0x0C51
        "10001011", -- 0x0C52
        "11100101", -- 0x0C53
        "10010011", -- 0x0C54
        "11111111", -- 0x0C55
        "10010000", -- 0x0C56
        "00000001", -- 0x0C57
        "00100011", -- 0x0C58
        "01111110", -- 0x0C59
        "00000000", -- 0x0C5A
        "00010010", -- 0x0C5B
        "00011111", -- 0x0C5C
        "10010001", -- 0x0C5D
        "10010000", -- 0x0C5E
        "00000001", -- 0x0C5F
        "00100011", -- 0x0C60
        "11100000", -- 0x0C61
        "11111110", -- 0x0C62
        "10100011", -- 0x0C63
        "11100000", -- 0x0C64
        "11111111", -- 0x0C65
        "00010010", -- 0x0C66
        "00100100", -- 0x0C67
        "10010101", -- 0x0C68
        "00010010", -- 0x0C69
        "00001110", -- 0x0C6A
        "10011100", -- 0x0C6B
        "10010000", -- 0x0C6C
        "00000001", -- 0x0C6D
        "00011010", -- 0x0C6E
        "11100000", -- 0x0C6F
        "01110000", -- 0x0C70
        "00000101", -- 0x0C71
        "00010010", -- 0x0C72
        "00011000", -- 0x0C73
        "10010001", -- 0x0C74
        "10000000", -- 0x0C75
        "10111000", -- 0x0C76
        "10010000", -- 0x0C77
        "00000001", -- 0x0C78
        "00011010", -- 0x0C79
        "11100000", -- 0x0C7A
        "11111000", -- 0x0C7B
        "10110100", -- 0x0C7C
        "00000110", -- 0x0C7D
        "00001111", -- 0x0C7E
        "11100101", -- 0x0C7F
        "11101101", -- 0x0C80
        "01010100", -- 0x0C81
        "11000000", -- 0x0C82
        "01100100", -- 0x0C83
        "01000000", -- 0x0C84
        "00100100", -- 0x0C85
        "11111111", -- 0x0C86
        "10110011", -- 0x0C87
        "11100100", -- 0x0C88
        "00110011", -- 0x0C89
        "01110000", -- 0x0C8A
        "10100011", -- 0x0C8B
        "10000000", -- 0x0C8C
        "00001110", -- 0x0C8D
        "10111000", -- 0x0C8E
        "00001001", -- 0x0C8F
        "10011110", -- 0x0C90
        "00010010", -- 0x0C91
        "00011001", -- 0x0C92
        "01001000", -- 0x0C93
        "10010000", -- 0x0C94
        "00000001", -- 0x0C95
        "00101101", -- 0x0C96
        "00010010", -- 0x0C97
        "00100011", -- 0x0C98
        "10101011", -- 0x0C99
        "01000000", -- 0x0C9A
        "10010011", -- 0x0C9B
        "10010000", -- 0x0C9C
        "00000001", -- 0x0C9D
        "00011010", -- 0x0C9E
        "11100100", -- 0x0C9F
        "11110000", -- 0x0CA0
        "10000000", -- 0x0CA1
        "10001100", -- 0x0CA2
        "00010010", -- 0x0CA3
        "00011001", -- 0x0CA4
        "01001000", -- 0x0CA5
        "10010000", -- 0x0CA6
        "00000001", -- 0x0CA7
        "10001001", -- 0x0CA8
        "00010010", -- 0x0CA9
        "00100001", -- 0x0CAA
        "11001000", -- 0x0CAB
        "00010010", -- 0x0CAC
        "00100100", -- 0x0CAD
        "01101001", -- 0x0CAE
        "10010000", -- 0x0CAF
        "00000001", -- 0x0CB0
        "10010101", -- 0x0CB1
        "11110000", -- 0x0CB2
        "01010011", -- 0x0CB3
        "11010101", -- 0x0CB4
        "11001111", -- 0x0CB5
        "01000011", -- 0x0CB6
        "11010101", -- 0x0CB7
        "00010000", -- 0x0CB8
        "01110101", -- 0x0CB9
        "11010100", -- 0x0CBA
        "00000001", -- 0x0CBB
        "00010010", -- 0x0CBC
        "00100000", -- 0x0CBD
        "01011001", -- 0x0CBE
        "10010000", -- 0x0CBF
        "00000001", -- 0x0CC0
        "10101111", -- 0x0CC1
        "00010010", -- 0x0CC2
        "00100100", -- 0x0CC3
        "01010100", -- 0x0CC4
        "10010000", -- 0x0CC5
        "00000001", -- 0x0CC6
        "10101111", -- 0x0CC7
        "00010010", -- 0x0CC8
        "00100010", -- 0x0CC9
        "10110101", -- 0x0CCA
        "10010000", -- 0x0CCB
        "00000001", -- 0x0CCC
        "10101111", -- 0x0CCD
        "01111110", -- 0x0CCE
        "00000000", -- 0x0CCF
        "00010010", -- 0x0CD0
        "00011111", -- 0x0CD1
        "10010001", -- 0x0CD2
        "01010011", -- 0x0CD3
        "11010101", -- 0x0CD4
        "11001111", -- 0x0CD5
        "01000011", -- 0x0CD6
        "11010101", -- 0x0CD7
        "00100000", -- 0x0CD8
        "01010011", -- 0x0CD9
        "11010101", -- 0x0CDA
        "11110011", -- 0x0CDB
        "01000011", -- 0x0CDC
        "11010101", -- 0x0CDD
        "00000100", -- 0x0CDE
        "01110101", -- 0x0CDF
        "11010100", -- 0x0CE0
        "00000011", -- 0x0CE1
        "00010010", -- 0x0CE2
        "00100000", -- 0x0CE3
        "01011001", -- 0x0CE4
        "10010000", -- 0x0CE5
        "00000001", -- 0x0CE6
        "10101101", -- 0x0CE7
        "00010010", -- 0x0CE8
        "00100100", -- 0x0CE9
        "01010100", -- 0x0CEA
        "10010000", -- 0x0CEB
        "00000001", -- 0x0CEC
        "10101101", -- 0x0CED
        "00010010", -- 0x0CEE
        "00100010", -- 0x0CEF
        "10110101", -- 0x0CF0
        "10010000", -- 0x0CF1
        "00000001", -- 0x0CF2
        "10101101", -- 0x0CF3
        "01111110", -- 0x0CF4
        "00000000", -- 0x0CF5
        "00010010", -- 0x0CF6
        "00011111", -- 0x0CF7
        "10010001", -- 0x0CF8
        "01010011", -- 0x0CF9
        "11010101", -- 0x0CFA
        "11110011", -- 0x0CFB
        "01000011", -- 0x0CFC
        "11010101", -- 0x0CFD
        "00001000", -- 0x0CFE
        "01110101", -- 0x0CFF
        "11010100", -- 0x0D00
        "00000000", -- 0x0D01
        "00010010", -- 0x0D02
        "00100100", -- 0x0D03
        "01101110", -- 0x0D04
        "10010000", -- 0x0D05
        "00000001", -- 0x0D06
        "10100010", -- 0x0D07
        "11110000", -- 0x0D08
        "01111110", -- 0x0D09
        "00010111", -- 0x0D0A
        "01111111", -- 0x0D0B
        "11111101", -- 0x0D0C
        "00010010", -- 0x0D0D
        "00010111", -- 0x0D0E
        "00000111", -- 0x0D0F
        "10010000", -- 0x0D10
        "00010111", -- 0x0D11
        "11111101", -- 0x0D12
        "11100000", -- 0x0D13
        "10010000", -- 0x0D14
        "00000001", -- 0x0D15
        "10100011", -- 0x0D16
        "11110000", -- 0x0D17
        "10010000", -- 0x0D18
        "00010111", -- 0x0D19
        "11111110", -- 0x0D1A
        "11100000", -- 0x0D1B
        "10010000", -- 0x0D1C
        "00000001", -- 0x0D1D
        "10100100", -- 0x0D1E
        "11110000", -- 0x0D1F
        "10010000", -- 0x0D20
        "00010111", -- 0x0D21
        "11111111", -- 0x0D22
        "00010010", -- 0x0D23
        "00100001", -- 0x0D24
        "10111100", -- 0x0D25
        "10010000", -- 0x0D26
        "00000001", -- 0x0D27
        "10100101", -- 0x0D28
        "00010010", -- 0x0D29
        "00100001", -- 0x0D2A
        "11001000", -- 0x0D2B
        "10010000", -- 0x0D2C
        "00011000", -- 0x0D2D
        "00000011", -- 0x0D2E
        "00010010", -- 0x0D2F
        "00100001", -- 0x0D30
        "10111100", -- 0x0D31
        "10010000", -- 0x0D32
        "00000001", -- 0x0D33
        "10101001", -- 0x0D34
        "00010010", -- 0x0D35
        "00100001", -- 0x0D36
        "11001000", -- 0x0D37
        "01111100", -- 0x0D38
        "00000000", -- 0x0D39
        "01111101", -- 0x0D3A
        "00101111", -- 0x0D3B
        "01111110", -- 0x0D3C
        "00000001", -- 0x0D3D
        "01111111", -- 0x0D3E
        "10000101", -- 0x0D3F
        "00010010", -- 0x0D40
        "00010111", -- 0x0D41
        "10001110", -- 0x0D42
        "10010000", -- 0x0D43
        "00000001", -- 0x0D44
        "10110100", -- 0x0D45
        "11110000", -- 0x0D46
        "00010010", -- 0x0D47
        "00100010", -- 0x0D48
        "00010111", -- 0x0D49
        "10010000", -- 0x0D4A
        "00000001", -- 0x0D4B
        "10000111", -- 0x0D4C
        "00010010", -- 0x0D4D
        "00011111", -- 0x0D4E
        "01011000", -- 0x0D4F
        "01110100", -- 0x0D50
        "11111111", -- 0x0D51
        "00100010", -- 0x0D52
        "10001111", -- 0x0D53
        "00001001", -- 0x0D54
        "10001110", -- 0x0D55
        "00001000", -- 0x0D56
        "01110101", -- 0x0D57
        "00001010", -- 0x0D58
        "00010101", -- 0x0D59
        "00010010", -- 0x0D5A
        "00100100", -- 0x0D5B
        "00100100", -- 0x0D5C
        "01100000", -- 0x0D5D
        "01111100", -- 0x0D5E
        "10000101", -- 0x0D5F
        "00001001", -- 0x0D60
        "10000010", -- 0x0D61
        "10000101", -- 0x0D62
        "00001000", -- 0x0D63
        "10000011", -- 0x0D64
        "11100000", -- 0x0D65
        "01100000", -- 0x0D66
        "00100010", -- 0x0D67
        "00100100", -- 0x0D68
        "11101011", -- 0x0D69
        "01100000", -- 0x0D6A
        "00110101", -- 0x0D6B
        "00100100", -- 0x0D6C
        "11110111", -- 0x0D6D
        "01100000", -- 0x0D6E
        "00101000", -- 0x0D6F
        "00100100", -- 0x0D70
        "11110001", -- 0x0D71
        "01100000", -- 0x0D72
        "01000010", -- 0x0D73
        "00100100", -- 0x0D74
        "11111010", -- 0x0D75
        "01100000", -- 0x0D76
        "01001100", -- 0x0D77
        "00100100", -- 0x0D78
        "11101000", -- 0x0D79
        "01100000", -- 0x0D7A
        "01010001", -- 0x0D7B
        "00100100", -- 0x0D7C
        "11000100", -- 0x0D7D
        "01100000", -- 0x0D7E
        "00001111", -- 0x0D7F
        "00100100", -- 0x0D80
        "11101110", -- 0x0D81
        "01100000", -- 0x0D82
        "00110111", -- 0x0D83
        "00100100", -- 0x0D84
        "11101111", -- 0x0D85
        "01100000", -- 0x0D86
        "00100101", -- 0x0D87
        "10000000", -- 0x0D88
        "01001100", -- 0x0D89
        "01110101", -- 0x0D8A
        "00001010", -- 0x0D8B
        "00000000", -- 0x0D8C
        "10000000", -- 0x0D8D
        "01000111", -- 0x0D8E
        "10101111", -- 0x0D8F
        "00001001", -- 0x0D90
        "10101110", -- 0x0D91
        "00001000", -- 0x0D92
        "00010010", -- 0x0D93
        "00011000", -- 0x0D94
        "00010010", -- 0x0D95
        "10000000", -- 0x0D96
        "00111100", -- 0x0D97
        "10101111", -- 0x0D98
        "00001001", -- 0x0D99
        "10101110", -- 0x0D9A
        "00001000", -- 0x0D9B
        "00010010", -- 0x0D9C
        "00000001", -- 0x0D9D
        "01001111", -- 0x0D9E
        "10000000", -- 0x0D9F
        "00110011", -- 0x0DA0
        "10101111", -- 0x0DA1
        "00001001", -- 0x0DA2
        "10101110", -- 0x0DA3
        "00001000", -- 0x0DA4
        "00010010", -- 0x0DA5
        "00000001", -- 0x0DA6
        "01001111", -- 0x0DA7
        "01110101", -- 0x0DA8
        "00001010", -- 0x0DA9
        "11111111", -- 0x0DAA
        "10000000", -- 0x0DAB
        "00101001", -- 0x0DAC
        "10101111", -- 0x0DAD
        "00001001", -- 0x0DAE
        "10101110", -- 0x0DAF
        "00001000", -- 0x0DB0
        "00010010", -- 0x0DB1
        "00010111", -- 0x0DB2
        "01001011", -- 0x0DB3
        "10000000", -- 0x0DB4
        "00011110", -- 0x0DB5
        "00010010", -- 0x0DB6
        "00001100", -- 0x0DB7
        "10100011", -- 0x0DB8
        "10000000", -- 0x0DB9
        "00011001", -- 0x0DBA
        "10101111", -- 0x0DBB
        "00001001", -- 0x0DBC
        "10101110", -- 0x0DBD
        "00001000", -- 0x0DBE
        "00010010", -- 0x0DBF
        "00000111", -- 0x0DC0
        "10001001", -- 0x0DC1
        "10000000", -- 0x0DC2
        "00010000", -- 0x0DC3
        "10101111", -- 0x0DC4
        "00001001", -- 0x0DC5
        "10101110", -- 0x0DC6
        "00001000", -- 0x0DC7
        "00010010", -- 0x0DC8
        "00011010", -- 0x0DC9
        "10111011", -- 0x0DCA
        "10000000", -- 0x0DCB
        "00000111", -- 0x0DCC
        "10101111", -- 0x0DCD
        "00001001", -- 0x0DCE
        "10101110", -- 0x0DCF
        "00001000", -- 0x0DD0
        "00010010", -- 0x0DD1
        "00010010", -- 0x0DD2
        "11011000", -- 0x0DD3
        "11110101", -- 0x0DD4
        "00001010", -- 0x0DD5
        "10101111", -- 0x0DD6
        "00001010", -- 0x0DD7
        "00000010", -- 0x0DD8
        "00011000", -- 0x0DD9
        "01010010", -- 0x0DDA
        "10000101", -- 0x0DDB
        "00001001", -- 0x0DDC
        "10000010", -- 0x0DDD
        "10000101", -- 0x0DDE
        "00001000", -- 0x0DDF
        "10000011", -- 0x0DE0
        "11100000", -- 0x0DE1
        "10110100", -- 0x0DE2
        "10000111", -- 0x0DE3
        "00000111", -- 0x0DE4
        "10101111", -- 0x0DE5
        "00001001", -- 0x0DE6
        "10101110", -- 0x0DE7
        "00001000", -- 0x0DE8
        "00000010", -- 0x0DE9
        "00011000", -- 0x0DEA
        "00010010", -- 0x0DEB
        "11100100", -- 0x0DEC
        "11111111", -- 0x0DED
        "11111110", -- 0x0DEE
        "11111101", -- 0x0DEF
        "11111100", -- 0x0DF0
        "00010010", -- 0x0DF1
        "00100100", -- 0x0DF2
        "00010010", -- 0x0DF3
        "01111111", -- 0x0DF4
        "01000000", -- 0x0DF5
        "00000010", -- 0x0DF6
        "00010001", -- 0x0DF7
        "11110101", -- 0x0DF8
        "10010000", -- 0x0DF9
        "00011000", -- 0x0DFA
        "00110001", -- 0x0DFB
        "00010010", -- 0x0DFC
        "00100001", -- 0x0DFD
        "01110100", -- 0x0DFE
        "10010000", -- 0x0DFF
        "00000000", -- 0x0E00
        "00000110", -- 0x0E01
        "11100000", -- 0x0E02
        "11111110", -- 0x0E03
        "10100011", -- 0x0E04
        "11100000", -- 0x0E05
        "11111111", -- 0x0E06
        "00010010", -- 0x0E07
        "00100100", -- 0x0E08
        "10010101", -- 0x0E09
        "10010000", -- 0x0E0A
        "00000001", -- 0x0E0B
        "00111001", -- 0x0E0C
        "00010010", -- 0x0E0D
        "00100001", -- 0x0E0E
        "11001000", -- 0x0E0F
        "11100100", -- 0x0E10
        "01111111", -- 0x0E11
        "11101000", -- 0x0E12
        "01111110", -- 0x0E13
        "00000011", -- 0x0E14
        "11111101", -- 0x0E15
        "11111100", -- 0x0E16
        "10010000", -- 0x0E17
        "00000001", -- 0x0E18
        "00111001", -- 0x0E19
        "00010010", -- 0x0E1A
        "00001001", -- 0x0E1B
        "10000110", -- 0x0E1C
        "10010000", -- 0x0E1D
        "00000001", -- 0x0E1E
        "00111001", -- 0x0E1F
        "00010010", -- 0x0E20
        "00100001", -- 0x0E21
        "11001000", -- 0x0E22
        "10010000", -- 0x0E23
        "00011000", -- 0x0E24
        "00110001", -- 0x0E25
        "00010010", -- 0x0E26
        "00100001", -- 0x0E27
        "10111100", -- 0x0E28
        "01110100", -- 0x0E29
        "00000001", -- 0x0E2A
        "00010010", -- 0x0E2B
        "00011111", -- 0x0E2C
        "00011100", -- 0x0E2D
        "10010000", -- 0x0E2E
        "00000001", -- 0x0E2F
        "00111001", -- 0x0E30
        "00010010", -- 0x0E31
        "00011011", -- 0x0E32
        "11010001", -- 0x0E33
        "10010000", -- 0x0E34
        "00011000", -- 0x0E35
        "00110001", -- 0x0E36
        "00010010", -- 0x0E37
        "00100001", -- 0x0E38
        "10111100", -- 0x0E39
        "10010000", -- 0x0E3A
        "00000001", -- 0x0E3B
        "00111001", -- 0x0E3C
        "00010010", -- 0x0E3D
        "00011010", -- 0x0E3E
        "01011110", -- 0x0E3F
        "10010000", -- 0x0E40
        "00000001", -- 0x0E41
        "00111001", -- 0x0E42
        "00010010", -- 0x0E43
        "00011011", -- 0x0E44
        "10000100", -- 0x0E45
        "10010000", -- 0x0E46
        "00000001", -- 0x0E47
        "00111001", -- 0x0E48
        "00010010", -- 0x0E49
        "00100001", -- 0x0E4A
        "10111100", -- 0x0E4B
        "10010000", -- 0x0E4C
        "00011000", -- 0x0E4D
        "00110101", -- 0x0E4E
        "00010010", -- 0x0E4F
        "00100001", -- 0x0E50
        "11001000", -- 0x0E51
        "10010000", -- 0x0E52
        "00000001", -- 0x0E53
        "00111001", -- 0x0E54
        "00010010", -- 0x0E55
        "00100001", -- 0x0E56
        "01010000", -- 0x0E57
        "10010000", -- 0x0E58
        "00000001", -- 0x0E59
        "00111100", -- 0x0E5A
        "11100000", -- 0x0E5B
        "11110101", -- 0x0E5C
        "11110111", -- 0x0E5D
        "01110101", -- 0x0E5E
        "10001001", -- 0x0E5F
        "01100110", -- 0x0E60
        "01110101", -- 0x0E61
        "10001000", -- 0x0E62
        "01010000", -- 0x0E63
        "01110101", -- 0x0E64
        "10001100", -- 0x0E65
        "11111111", -- 0x0E66
        "01110101", -- 0x0E67
        "10001101", -- 0x0E68
        "11111111", -- 0x0E69
        "01110101", -- 0x0E6A
        "10001010", -- 0x0E6B
        "11111111", -- 0x0E6C
        "01110101", -- 0x0E6D
        "10001011", -- 0x0E6E
        "11111111", -- 0x0E6F
        "11000010", -- 0x0E70
        "10111001", -- 0x0E71
        "11010010", -- 0x0E72
        "10101011", -- 0x0E73
        "11000010", -- 0x0E74
        "10101001", -- 0x0E75
        "11010010", -- 0x0E76
        "10101000", -- 0x0E77
        "11010010", -- 0x0E78
        "10001000", -- 0x0E79
        "11010010", -- 0x0E7A
        "10101010", -- 0x0E7B
        "11010010", -- 0x0E7C
        "10001010", -- 0x0E7D
        "11010010", -- 0x0E7E
        "10111010", -- 0x0E7F
        "11010010", -- 0x0E80
        "10101111", -- 0x0E81
        "11100100", -- 0x0E82
        "01111111", -- 0x0E83
        "00000001", -- 0x0E84
        "11111110", -- 0x0E85
        "11111101", -- 0x0E86
        "11111100", -- 0x0E87
        "00010010", -- 0x0E88
        "00010110", -- 0x0E89
        "00110100", -- 0x0E8A
        "10010000", -- 0x0E8B
        "00000000", -- 0x0E8C
        "00000001", -- 0x0E8D
        "01110100", -- 0x0E8E
        "00000001", -- 0x0E8F
        "11110000", -- 0x0E90
        "10010000", -- 0x0E91
        "00000000", -- 0x0E92
        "00000000", -- 0x0E93
        "00010100", -- 0x0E94
        "11110000", -- 0x0E95
        "10010000", -- 0x0E96
        "00000000", -- 0x0E97
        "00000010", -- 0x0E98
        "11100100", -- 0x0E99
        "11110000", -- 0x0E9A
        "00100010", -- 0x0E9B
        "10010000", -- 0x0E9C
        "00011000", -- 0x0E9D
        "00101001", -- 0x0E9E
        "00010010", -- 0x0E9F
        "00100001", -- 0x0EA0
        "01110100", -- 0x0EA1
        "11100100", -- 0x0EA2
        "11111110", -- 0x0EA3
        "11111101", -- 0x0EA4
        "11111100", -- 0x0EA5
        "10010000", -- 0x0EA6
        "00011000", -- 0x0EA7
        "00101001", -- 0x0EA8
        "01111111", -- 0x0EA9
        "01100000", -- 0x0EAA
        "00010010", -- 0x0EAB
        "00001001", -- 0x0EAC
        "10000110", -- 0x0EAD
        "10010000", -- 0x0EAE
        "00011000", -- 0x0EAF
        "00101101", -- 0x0EB0
        "00010010", -- 0x0EB1
        "00100001", -- 0x0EB2
        "11001000", -- 0x0EB3
        "00010010", -- 0x0EB4
        "00100010", -- 0x0EB5
        "10000110", -- 0x0EB6
        "00010010", -- 0x0EB7
        "00011101", -- 0x0EB8
        "11000011", -- 0x0EB9
        "10101001", -- 0x0EBA
        "00000111", -- 0x0EBB
        "10101000", -- 0x0EBC
        "00000110", -- 0x0EBD
        "00010010", -- 0x0EBE
        "00100010", -- 0x0EBF
        "10000110", -- 0x0EC0
        "00010010", -- 0x0EC1
        "00011101", -- 0x0EC2
        "11011110", -- 0x0EC3
        "11101111", -- 0x0EC4
        "00100100", -- 0x0EC5
        "11111010", -- 0x0EC6
        "11101110", -- 0x0EC7
        "00110100", -- 0x0EC8
        "11111111", -- 0x0EC9
        "11101101", -- 0x0ECA
        "00110100", -- 0x0ECB
        "11111111", -- 0x0ECC
        "11101100", -- 0x0ECD
        "00110100", -- 0x0ECE
        "11111111", -- 0x0ECF
        "01010000", -- 0x0ED0
        "00000100", -- 0x0ED1
        "01110100", -- 0x0ED2
        "00000001", -- 0x0ED3
        "10000000", -- 0x0ED4
        "00000001", -- 0x0ED5
        "11100100", -- 0x0ED6
        "11111011", -- 0x0ED7
        "01111010", -- 0x0ED8
        "00000000", -- 0x0ED9
        "11101001", -- 0x0EDA
        "00101011", -- 0x0EDB
        "11111001", -- 0x0EDC
        "11101000", -- 0x0EDD
        "00111010", -- 0x0EDE
        "11111000", -- 0x0EDF
        "11110101", -- 0x0EE0
        "10100011", -- 0x0EE1
        "11101001", -- 0x0EE2
        "11110101", -- 0x0EE3
        "10101011", -- 0x0EE4
        "10001001", -- 0x0EE5
        "00000111", -- 0x0EE6
        "10001000", -- 0x0EE7
        "00000110", -- 0x0EE8
        "00010010", -- 0x0EE9
        "00100100", -- 0x0EEA
        "10010101", -- 0x0EEB
        "00010010", -- 0x0EEC
        "00100001", -- 0x0EED
        "00011110", -- 0x0EEE
        "01111110", -- 0x0EEF
        "00000011", -- 0x0EF0
        "01111111", -- 0x0EF1
        "11101000", -- 0x0EF2
        "00010010", -- 0x0EF3
        "00001001", -- 0x0EF4
        "10000110", -- 0x0EF5
        "00010010", -- 0x0EF6
        "00100001", -- 0x0EF7
        "00011110", -- 0x0EF8
        "01111110", -- 0x0EF9
        "00010010", -- 0x0EFA
        "01111111", -- 0x0EFB
        "11000000", -- 0x0EFC
        "00010010", -- 0x0EFD
        "00011011", -- 0x0EFE
        "11010001", -- 0x0EFF
        "11100100", -- 0x0F00
        "11111101", -- 0x0F01
        "11111100", -- 0x0F02
        "10010000", -- 0x0F03
        "00011000", -- 0x0F04
        "00101101", -- 0x0F05
        "01111110", -- 0x0F06
        "00100101", -- 0x0F07
        "01111111", -- 0x0F08
        "10000000", -- 0x0F09
        "00010010", -- 0x0F0A
        "00011010", -- 0x0F0B
        "01011110", -- 0x0F0C
        "10010000", -- 0x0F0D
        "00011000", -- 0x0F0E
        "00101101", -- 0x0F0F
        "00010010", -- 0x0F10
        "00011011", -- 0x0F11
        "10000100", -- 0x0F12
        "10010000", -- 0x0F13
        "00011000", -- 0x0F14
        "00101101", -- 0x0F15
        "00010010", -- 0x0F16
        "00100001", -- 0x0F17
        "01010000", -- 0x0F18
        "10010000", -- 0x0F19
        "00011000", -- 0x0F1A
        "00110000", -- 0x0F1B
        "11100000", -- 0x0F1C
        "11110101", -- 0x0F1D
        "11110111", -- 0x0F1E
        "01000011", -- 0x0F1F
        "11001100", -- 0x0F20
        "00000010", -- 0x0F21
        "01010011", -- 0x0F22
        "11001100", -- 0x0F23
        "11111101", -- 0x0F24
        "10010000", -- 0x0F25
        "00000000", -- 0x0F26
        "00000110", -- 0x0F27
        "11101000", -- 0x0F28
        "11110000", -- 0x0F29
        "11101001", -- 0x0F2A
        "10100011", -- 0x0F2B
        "11110000", -- 0x0F2C
        "10010000", -- 0x0F2D
        "00011000", -- 0x0F2E
        "00101101", -- 0x0F2F
        "00010010", -- 0x0F30
        "00100001", -- 0x0F31
        "10111100", -- 0x0F32
        "10010000", -- 0x0F33
        "00000001", -- 0x0F34
        "00110101", -- 0x0F35
        "00000010", -- 0x0F36
        "00100001", -- 0x0F37
        "11001000", -- 0x0F38
        "10010000", -- 0x0F39
        "00000001", -- 0x0F3A
        "00011011", -- 0x0F3B
        "11100000", -- 0x0F3C
        "01100000", -- 0x0F3D
        "00000011", -- 0x0F3E
        "00000010", -- 0x0F3F
        "00001111", -- 0x0F40
        "11010011", -- 0x0F41
        "10010000", -- 0x0F42
        "00000000", -- 0x0F43
        "00010000", -- 0x0F44
        "11100000", -- 0x0F45
        "01110000", -- 0x0F46
        "00011101", -- 0x0F47
        "10010000", -- 0x0F48
        "00000000", -- 0x0F49
        "00010001", -- 0x0F4A
        "11100000", -- 0x0F4B
        "10110100", -- 0x0F4C
        "11111111", -- 0x0F4D
        "00010110", -- 0x0F4E
        "01111001", -- 0x0F4F
        "00010000", -- 0x0F50
        "01111000", -- 0x0F51
        "00000000", -- 0x0F52
        "01111010", -- 0x0F53
        "00001000", -- 0x0F54
        "10010000", -- 0x0F55
        "00000001", -- 0x0F56
        "10010110", -- 0x0F57
        "11100000", -- 0x0F58
        "10001001", -- 0x0F59
        "10000010", -- 0x0F5A
        "10001000", -- 0x0F5B
        "10000011", -- 0x0F5C
        "11110000", -- 0x0F5D
        "00001001", -- 0x0F5E
        "10111001", -- 0x0F5F
        "00000000", -- 0x0F60
        "00000001", -- 0x0F61
        "00001000", -- 0x0F62
        "11011010", -- 0x0F63
        "11110000", -- 0x0F64
        "01111001", -- 0x0F65
        "00010001", -- 0x0F66
        "01111000", -- 0x0F67
        "00000000", -- 0x0F68
        "01111011", -- 0x0F69
        "00010000", -- 0x0F6A
        "01111010", -- 0x0F6B
        "00000000", -- 0x0F6C
        "01111100", -- 0x0F6D
        "00000111", -- 0x0F6E
        "10001001", -- 0x0F6F
        "10000010", -- 0x0F70
        "10001000", -- 0x0F71
        "10000011", -- 0x0F72
        "11100000", -- 0x0F73
        "10001011", -- 0x0F74
        "10000010", -- 0x0F75
        "10001010", -- 0x0F76
        "10000011", -- 0x0F77
        "11110000", -- 0x0F78
        "00001011", -- 0x0F79
        "10111011", -- 0x0F7A
        "00000000", -- 0x0F7B
        "00000001", -- 0x0F7C
        "00001010", -- 0x0F7D
        "00001001", -- 0x0F7E
        "10111001", -- 0x0F7F
        "00000000", -- 0x0F80
        "00000001", -- 0x0F81
        "00001000", -- 0x0F82
        "11011100", -- 0x0F83
        "11101010", -- 0x0F84
        "10010000", -- 0x0F85
        "00000001", -- 0x0F86
        "10010110", -- 0x0F87
        "11100000", -- 0x0F88
        "10010000", -- 0x0F89
        "00000000", -- 0x0F8A
        "00010111", -- 0x0F8B
        "11110000", -- 0x0F8C
        "10010000", -- 0x0F8D
        "00000000", -- 0x0F8E
        "00010000", -- 0x0F8F
        "00010010", -- 0x0F90
        "00011111", -- 0x0F91
        "11000110", -- 0x0F92
        "10010000", -- 0x0F93
        "00000000", -- 0x0F94
        "00010011", -- 0x0F95
        "00010010", -- 0x0F96
        "00100001", -- 0x0F97
        "10000000", -- 0x0F98
        "10001111", -- 0x0F99
        "00010011", -- 0x0F9A
        "10001110", -- 0x0F9B
        "00010010", -- 0x0F9C
        "10010000", -- 0x0F9D
        "00000000", -- 0x0F9E
        "00010100", -- 0x0F9F
        "00010010", -- 0x0FA0
        "00011111", -- 0x0FA1
        "11000110", -- 0x0FA2
        "10010000", -- 0x0FA3
        "00000000", -- 0x0FA4
        "00010111", -- 0x0FA5
        "00010010", -- 0x0FA6
        "00100001", -- 0x0FA7
        "10000000", -- 0x0FA8
        "11100101", -- 0x0FA9
        "00010011", -- 0x0FAA
        "11010011", -- 0x0FAB
        "10011111", -- 0x0FAC
        "11100101", -- 0x0FAD
        "00010010", -- 0x0FAE
        "10011110", -- 0x0FAF
        "01000000", -- 0x0FB0
        "00100001", -- 0x0FB1
        "11100101", -- 0x0FB2
        "00010011", -- 0x0FB3
        "11000011", -- 0x0FB4
        "10011111", -- 0x0FB5
        "11111001", -- 0x0FB6
        "11100101", -- 0x0FB7
        "00010010", -- 0x0FB8
        "10011110", -- 0x0FB9
        "11111000", -- 0x0FBA
        "11101001", -- 0x0FBB
        "00100100", -- 0x0FBC
        "11111110", -- 0x0FBD
        "11101000", -- 0x0FBE
        "00110100", -- 0x0FBF
        "11111111", -- 0x0FC0
        "01010000", -- 0x0FC1
        "00010000", -- 0x0FC2
        "10010000", -- 0x0FC3
        "00000001", -- 0x0FC4
        "00011011", -- 0x0FC5
        "01110100", -- 0x0FC6
        "00000001", -- 0x0FC7
        "11110000", -- 0x0FC8
        "11100100", -- 0x0FC9
        "11111101", -- 0x0FCA
        "11111100", -- 0x0FCB
        "01111110", -- 0x0FCC
        "00001111", -- 0x0FCD
        "01111111", -- 0x0FCE
        "00111001", -- 0x0FCF
        "00010010", -- 0x0FD0
        "00010100", -- 0x0FD1
        "00010100", -- 0x0FD2
        "00100010", -- 0x0FD3
        "10111100", -- 0x0FD4
        "00000000", -- 0x0FD5
        "00010100", -- 0x0FD6
        "10111101", -- 0x0FD7
        "00000000", -- 0x0FD8
        "00000010", -- 0x0FD9
        "11010011", -- 0x0FDA
        "00100010", -- 0x0FDB
        "10111110", -- 0x0FDC
        "00000000", -- 0x0FDD
        "01001111", -- 0x0FDE
        "11000101", -- 0x0FDF
        "11110000", -- 0x0FE0
        "10001101", -- 0x0FE1
        "11110000", -- 0x0FE2
        "11001111", -- 0x0FE3
        "10000100", -- 0x0FE4
        "11001111", -- 0x0FE5
        "10101101", -- 0x0FE6
        "11110000", -- 0x0FE7
        "11000101", -- 0x0FE8
        "11110000", -- 0x0FE9
        "00100010", -- 0x0FEA
        "10111110", -- 0x0FEB
        "00000000", -- 0x0FEC
        "00001000", -- 0x0FED
        "11101111", -- 0x0FEE
        "11111101", -- 0x0FEF
        "11101110", -- 0x0FF0
        "11111100", -- 0x0FF1
        "11100100", -- 0x0FF2
        "11111111", -- 0x0FF3
        "11111110", -- 0x0FF4
        "00100010", -- 0x0FF5
        "11000011", -- 0x0FF6
        "11101111", -- 0x0FF7
        "10011101", -- 0x0FF8
        "11101110", -- 0x0FF9
        "10011100", -- 0x0FFA
        "01000000", -- 0x0FFB
        "11110001", -- 0x0FFC
        "11000000", -- 0x0FFD
        "11110000", -- 0x0FFE
        "11101000", -- 0x0FFF
        "11000000", -- 0x1000
        "11100000", -- 0x1001
        "11101001", -- 0x1002
        "11000000", -- 0x1003
        "11100000", -- 0x1004
        "11100100", -- 0x1005
        "11111001", -- 0x1006
        "01111000", -- 0x1007
        "00000001", -- 0x1008
        "11000011", -- 0x1009
        "11101111", -- 0x100A
        "00110011", -- 0x100B
        "11111111", -- 0x100C
        "11101110", -- 0x100D
        "00110011", -- 0x100E
        "11111110", -- 0x100F
        "11101001", -- 0x1010
        "00110011", -- 0x1011
        "11111001", -- 0x1012
        "11101110", -- 0x1013
        "10011101", -- 0x1014
        "11110101", -- 0x1015
        "11110000", -- 0x1016
        "11101001", -- 0x1017
        "10011100", -- 0x1018
        "10110011", -- 0x1019
        "01010000", -- 0x101A
        "00000011", -- 0x101B
        "11111001", -- 0x101C
        "10101110", -- 0x101D
        "11110000", -- 0x101E
        "11101000", -- 0x101F
        "00110011", -- 0x1020
        "11111000", -- 0x1021
        "01010000", -- 0x1022
        "11100101", -- 0x1023
        "11101001", -- 0x1024
        "11111100", -- 0x1025
        "11101110", -- 0x1026
        "11111101", -- 0x1027
        "11101000", -- 0x1028
        "11111111", -- 0x1029
        "01111110", -- 0x102A
        "00000000", -- 0x102B
        "10000000", -- 0x102C
        "00110011", -- 0x102D
        "11000000", -- 0x102E
        "11110000", -- 0x102F
        "11101000", -- 0x1030
        "11000000", -- 0x1031
        "11100000", -- 0x1032
        "11101001", -- 0x1033
        "11000000", -- 0x1034
        "11100000", -- 0x1035
        "01111000", -- 0x1036
        "00001001", -- 0x1037
        "11101111", -- 0x1038
        "11111001", -- 0x1039
        "01111111", -- 0x103A
        "00000000", -- 0x103B
        "10001101", -- 0x103C
        "11110000", -- 0x103D
        "10101100", -- 0x103E
        "11110000", -- 0x103F
        "11101110", -- 0x1040
        "10000100", -- 0x1041
        "11111110", -- 0x1042
        "11100101", -- 0x1043
        "11110000", -- 0x1044
        "11000011", -- 0x1045
        "01010000", -- 0x1046
        "00000110", -- 0x1047
        "11001111", -- 0x1048
        "00110011", -- 0x1049
        "11001111", -- 0x104A
        "10011100", -- 0x104B
        "10000000", -- 0x104C
        "00001000", -- 0x104D
        "10011100", -- 0x104E
        "01010000", -- 0x104F
        "00000001", -- 0x1050
        "00101100", -- 0x1051
        "11001111", -- 0x1052
        "10110011", -- 0x1053
        "00110011", -- 0x1054
        "11001111", -- 0x1055
        "11001001", -- 0x1056
        "00100101", -- 0x1057
        "11100000", -- 0x1058
        "11001001", -- 0x1059
        "11111101", -- 0x105A
        "00110101", -- 0x105B
        "11100000", -- 0x105C
        "11011000", -- 0x105D
        "11100111", -- 0x105E
        "01111100", -- 0x105F
        "00000000", -- 0x1060
        "11010000", -- 0x1061
        "11100000", -- 0x1062
        "11111001", -- 0x1063
        "11010000", -- 0x1064
        "11100000", -- 0x1065
        "11111000", -- 0x1066
        "11010000", -- 0x1067
        "11110000", -- 0x1068
        "11000011", -- 0x1069
        "00100010", -- 0x106A
        "11101111", -- 0x106B
        "01001110", -- 0x106C
        "01001101", -- 0x106D
        "01001100", -- 0x106E
        "01110000", -- 0x106F
        "00000010", -- 0x1070
        "11010011", -- 0x1071
        "00100010", -- 0x1072
        "11101000", -- 0x1073
        "11000000", -- 0x1074
        "11100000", -- 0x1075
        "11101001", -- 0x1076
        "11000000", -- 0x1077
        "11100000", -- 0x1078
        "11101010", -- 0x1079
        "11000000", -- 0x107A
        "11100000", -- 0x107B
        "11101011", -- 0x107C
        "11000000", -- 0x107D
        "11100000", -- 0x107E
        "11100100", -- 0x107F
        "11000000", -- 0x1080
        "11100000", -- 0x1081
        "11000000", -- 0x1082
        "11100000", -- 0x1083
        "11000000", -- 0x1084
        "11100000", -- 0x1085
        "11000000", -- 0x1086
        "11100000", -- 0x1087
        "01111010", -- 0x1088
        "00100000", -- 0x1089
        "01111011", -- 0x108A
        "00000100", -- 0x108B
        "11100101", -- 0x108C
        "10000001", -- 0x108D
        "00100100", -- 0x108E
        "11110011", -- 0x108F
        "11111000", -- 0x1090
        "11100110", -- 0x1091
        "01110000", -- 0x1092
        "00010011", -- 0x1093
        "11101010", -- 0x1094
        "00100100", -- 0x1095
        "11111000", -- 0x1096
        "11111010", -- 0x1097
        "00001000", -- 0x1098
        "00001000", -- 0x1099
        "00001000", -- 0x109A
        "11100100", -- 0x109B
        "11000110", -- 0x109C
        "00011000", -- 0x109D
        "11000110", -- 0x109E
        "00011000", -- 0x109F
        "11000110", -- 0x10A0
        "00011000", -- 0x10A1
        "11110110", -- 0x10A2
        "11011011", -- 0x10A3
        "11101101", -- 0x10A4
        "10000000", -- 0x10A5
        "01000010", -- 0x10A6
        "01111011", -- 0x10A7
        "00000100", -- 0x10A8
        "11100101", -- 0x10A9
        "10000001", -- 0x10AA
        "11111001", -- 0x10AB
        "00100100", -- 0x10AC
        "11110110", -- 0x10AD
        "11111000", -- 0x10AE
        "11000011", -- 0x10AF
        "11100110", -- 0x10B0
        "00110011", -- 0x10B1
        "11110110", -- 0x10B2
        "00011000", -- 0x10B3
        "11011011", -- 0x10B4
        "11111010", -- 0x10B5
        "01111011", -- 0x10B6
        "00000100", -- 0x10B7
        "11100111", -- 0x10B8
        "00110011", -- 0x10B9
        "11110111", -- 0x10BA
        "00011001", -- 0x10BB
        "11011011", -- 0x10BC
        "11111010", -- 0x10BD
        "11000011", -- 0x10BE
        "11100101", -- 0x10BF
        "10000001", -- 0x10C0
        "11111000", -- 0x10C1
        "11100110", -- 0x10C2
        "10011111", -- 0x10C3
        "00011000", -- 0x10C4
        "11100110", -- 0x10C5
        "10011110", -- 0x10C6
        "00011000", -- 0x10C7
        "11100110", -- 0x10C8
        "10011101", -- 0x10C9
        "00011000", -- 0x10CA
        "11100110", -- 0x10CB
        "10011100", -- 0x10CC
        "01000000", -- 0x10CD
        "00011000", -- 0x10CE
        "11100101", -- 0x10CF
        "10000001", -- 0x10D0
        "00100100", -- 0x10D1
        "11110110", -- 0x10D2
        "11111000", -- 0x10D3
        "00000110", -- 0x10D4
        "11000011", -- 0x10D5
        "10101000", -- 0x10D6
        "10000001", -- 0x10D7
        "11100110", -- 0x10D8
        "10011111", -- 0x10D9
        "11110110", -- 0x10DA
        "00011000", -- 0x10DB
        "11100110", -- 0x10DC
        "10011110", -- 0x10DD
        "11110110", -- 0x10DE
        "00011000", -- 0x10DF
        "11100110", -- 0x10E0
        "10011101", -- 0x10E1
        "11110110", -- 0x10E2
        "00011000", -- 0x10E3
        "11100110", -- 0x10E4
        "10011100", -- 0x10E5
        "11110110", -- 0x10E6
        "11011010", -- 0x10E7
        "10111110", -- 0x10E8
        "11010000", -- 0x10E9
        "11100000", -- 0x10EA
        "11111111", -- 0x10EB
        "11010000", -- 0x10EC
        "11100000", -- 0x10ED
        "11111110", -- 0x10EE
        "11010000", -- 0x10EF
        "11100000", -- 0x10F0
        "11111101", -- 0x10F1
        "11010000", -- 0x10F2
        "11100000", -- 0x10F3
        "11111100", -- 0x10F4
        "11010000", -- 0x10F5
        "11100000", -- 0x10F6
        "11111011", -- 0x10F7
        "11010000", -- 0x10F8
        "11100000", -- 0x10F9
        "11111010", -- 0x10FA
        "11010000", -- 0x10FB
        "11100000", -- 0x10FC
        "11111001", -- 0x10FD
        "11010000", -- 0x10FE
        "11100000", -- 0x10FF
        "11111000", -- 0x1100
        "00100010", -- 0x1101
        "10001111", -- 0x1102
        "00000011", -- 0x1103
        "10001110", -- 0x1104
        "00000010", -- 0x1105
        "10001101", -- 0x1106
        "00011001", -- 0x1107
        "10001100", -- 0x1108
        "00011000", -- 0x1109
        "00010010", -- 0x110A
        "00100001", -- 0x110B
        "10011000", -- 0x110C
        "01110101", -- 0x110D
        "00010110", -- 0x110E
        "00000001", -- 0x110F
        "01110101", -- 0x1110
        "00010111", -- 0x1111
        "10110110", -- 0x1112
        "11100101", -- 0x1113
        "00010111", -- 0x1114
        "00101111", -- 0x1115
        "11111001", -- 0x1116
        "11100101", -- 0x1117
        "00010110", -- 0x1118
        "00111110", -- 0x1119
        "11111000", -- 0x111A
        "11101001", -- 0x111B
        "00100100", -- 0x111C
        "00000010", -- 0x111D
        "00010010", -- 0x111E
        "00100011", -- 0x111F
        "11101010", -- 0x1120
        "11100101", -- 0x1121
        "00011000", -- 0x1122
        "11110000", -- 0x1123
        "11100101", -- 0x1124
        "00011001", -- 0x1125
        "10100011", -- 0x1126
        "11110000", -- 0x1127
        "00010010", -- 0x1128
        "00100001", -- 0x1129
        "10110000", -- 0x112A
        "00010010", -- 0x112B
        "00100100", -- 0x112C
        "10000010", -- 0x112D
        "11101010", -- 0x112E
        "11110000", -- 0x112F
        "11101011", -- 0x1130
        "10100011", -- 0x1131
        "11110000", -- 0x1132
        "11100101", -- 0x1133
        "00011000", -- 0x1134
        "01000101", -- 0x1135
        "00011001", -- 0x1136
        "01100000", -- 0x1137
        "00101111", -- 0x1138
        "10101111", -- 0x1139
        "00011001", -- 0x113A
        "10101110", -- 0x113B
        "00011000", -- 0x113C
        "00010010", -- 0x113D
        "00000000", -- 0x113E
        "00000110", -- 0x113F
        "10001111", -- 0x1140
        "00000011", -- 0x1141
        "10001110", -- 0x1142
        "00000010", -- 0x1143
        "10001101", -- 0x1144
        "00000001", -- 0x1145
        "10001100", -- 0x1146
        "00000000", -- 0x1147
        "00010010", -- 0x1148
        "00100001", -- 0x1149
        "10011000", -- 0x114A
        "11100101", -- 0x114B
        "00010111", -- 0x114C
        "00101111", -- 0x114D
        "11111101", -- 0x114E
        "11100101", -- 0x114F
        "00010110", -- 0x1150
        "00111110", -- 0x1151
        "11111100", -- 0x1152
        "11101101", -- 0x1153
        "00100100", -- 0x1154
        "00000100", -- 0x1155
        "11111101", -- 0x1156
        "11100100", -- 0x1157
        "00111100", -- 0x1158
        "11111100", -- 0x1159
        "10001101", -- 0x115A
        "10000010", -- 0x115B
        "10001100", -- 0x115C
        "10000011", -- 0x115D
        "10001011", -- 0x115E
        "00000111", -- 0x115F
        "10001010", -- 0x1160
        "00000110", -- 0x1161
        "10001001", -- 0x1162
        "00000101", -- 0x1163
        "10001000", -- 0x1164
        "00000100", -- 0x1165
        "10000000", -- 0x1166
        "00001110", -- 0x1167
        "00010010", -- 0x1168
        "00100001", -- 0x1169
        "10110000", -- 0x116A
        "11101001", -- 0x116B
        "00100100", -- 0x116C
        "00000100", -- 0x116D
        "00010010", -- 0x116E
        "00100011", -- 0x116F
        "11101010", -- 0x1170
        "11100100", -- 0x1171
        "11111111", -- 0x1172
        "11111110", -- 0x1173
        "11111101", -- 0x1174
        "11111100", -- 0x1175
        "00010010", -- 0x1176
        "00100001", -- 0x1177
        "11001000", -- 0x1178
        "10010000", -- 0x1179
        "00000001", -- 0x117A
        "10110101", -- 0x117B
        "11100000", -- 0x117C
        "00000100", -- 0x117D
        "11110000", -- 0x117E
        "00100010", -- 0x117F
        "11000000", -- 0x1180
        "00000111", -- 0x1181
        "11000000", -- 0x1182
        "11100000", -- 0x1183
        "11000000", -- 0x1184
        "11110000", -- 0x1185
        "11000000", -- 0x1186
        "10000010", -- 0x1187
        "11000000", -- 0x1188
        "10000011", -- 0x1189
        "11000000", -- 0x118A
        "00000000", -- 0x118B
        "11000000", -- 0x118C
        "00000001", -- 0x118D
        "11000000", -- 0x118E
        "00000010", -- 0x118F
        "11000000", -- 0x1190
        "00000011", -- 0x1191
        "11000000", -- 0x1192
        "00000100", -- 0x1193
        "11000000", -- 0x1194
        "00000101", -- 0x1195
        "11000000", -- 0x1196
        "00000110", -- 0x1197
        "11000000", -- 0x1198
        "11010000", -- 0x1199
        "01110101", -- 0x119A
        "11010000", -- 0x119B
        "00000000", -- 0x119C
        "10010000", -- 0x119D
        "00000001", -- 0x119E
        "10010011", -- 0x119F
        "00010010", -- 0x11A0
        "00011111", -- 0x11A1
        "01011000", -- 0x11A2
        "10010000", -- 0x11A3
        "00000100", -- 0x11A4
        "10000100", -- 0x11A5
        "11100000", -- 0x11A6
        "10110100", -- 0x11A7
        "00000001", -- 0x11A8
        "00011111", -- 0x11A9
        "00010010", -- 0x11AA
        "00011001", -- 0x11AB
        "01001000", -- 0x11AC
        "10010000", -- 0x11AD
        "00000000", -- 0x11AE
        "00001000", -- 0x11AF
        "00010010", -- 0x11B0
        "00011010", -- 0x11B1
        "11100100", -- 0x11B2
        "10010000", -- 0x11B3
        "00011000", -- 0x11B4
        "00011100", -- 0x11B5
        "00010010", -- 0x11B6
        "00100001", -- 0x11B7
        "11001000", -- 0x11B8
        "10010000", -- 0x11B9
        "00011000", -- 0x11BA
        "00011110", -- 0x11BB
        "11100000", -- 0x11BC
        "11111000", -- 0x11BD
        "10100011", -- 0x11BE
        "11100000", -- 0x11BF
        "11111001", -- 0x11C0
        "10010000", -- 0x11C1
        "00000011", -- 0x11C2
        "10010010", -- 0x11C3
        "11101000", -- 0x11C4
        "11110000", -- 0x11C5
        "11101001", -- 0x11C6
        "10100011", -- 0x11C7
        "11110000", -- 0x11C8
        "10010000", -- 0x11C9
        "00000001", -- 0x11CA
        "10010110", -- 0x11CB
        "11100000", -- 0x11CC
        "11111111", -- 0x11CD
        "00010010", -- 0x11CE
        "00011001", -- 0x11CF
        "10000001", -- 0x11D0
        "00010010", -- 0x11D1
        "00011001", -- 0x11D2
        "01001000", -- 0x11D3
        "10010000", -- 0x11D4
        "00000000", -- 0x11D5
        "00001000", -- 0x11D6
        "00010010", -- 0x11D7
        "00100001", -- 0x11D8
        "11001000", -- 0x11D9
        "11010000", -- 0x11DA
        "11010000", -- 0x11DB
        "11010000", -- 0x11DC
        "00000110", -- 0x11DD
        "11010000", -- 0x11DE
        "00000101", -- 0x11DF
        "11010000", -- 0x11E0
        "00000100", -- 0x11E1
        "11010000", -- 0x11E2
        "00000011", -- 0x11E3
        "11010000", -- 0x11E4
        "00000010", -- 0x11E5
        "11010000", -- 0x11E6
        "00000001", -- 0x11E7
        "11010000", -- 0x11E8
        "00000000", -- 0x11E9
        "11010000", -- 0x11EA
        "10000011", -- 0x11EB
        "11010000", -- 0x11EC
        "10000010", -- 0x11ED
        "11010000", -- 0x11EE
        "11110000", -- 0x11EF
        "11010000", -- 0x11F0
        "11100000", -- 0x11F1
        "11010000", -- 0x11F2
        "00000111", -- 0x11F3
        "00110010", -- 0x11F4
        "10001111", -- 0x11F5
        "00001111", -- 0x11F6
        "00010010", -- 0x11F7
        "00011101", -- 0x11F8
        "10100111", -- 0x11F9
        "11100101", -- 0x11FA
        "00001111", -- 0x11FB
        "11110000", -- 0x11FC
        "10010000", -- 0x11FD
        "00010111", -- 0x11FE
        "11101001", -- 0x11FF
        "00010010", -- 0x1200
        "00100001", -- 0x1201
        "10111100", -- 0x1202
        "10010000", -- 0x1203
        "00010111", -- 0x1204
        "11100101", -- 0x1205
        "00010010", -- 0x1206
        "00100001", -- 0x1207
        "11001000", -- 0x1208
        "10010000", -- 0x1209
        "00000111", -- 0x120A
        "11001011", -- 0x120B
        "00010010", -- 0x120C
        "00011111", -- 0x120D
        "01011000", -- 0x120E
        "10010000", -- 0x120F
        "00000110", -- 0x1210
        "10001001", -- 0x1211
        "11100000", -- 0x1212
        "10110100", -- 0x1213
        "00100000", -- 0x1214
        "00111010", -- 0x1215
        "00010010", -- 0x1216
        "00100000", -- 0x1217
        "01001001", -- 0x1218
        "01110101", -- 0x1219
        "00001111", -- 0x121A
        "00000110", -- 0x121B
        "01110101", -- 0x121C
        "00010000", -- 0x121D
        "10001011", -- 0x121E
        "00100101", -- 0x121F
        "00010000", -- 0x1220
        "11111001", -- 0x1221
        "11101110", -- 0x1222
        "00110101", -- 0x1223
        "00001111", -- 0x1224
        "00010010", -- 0x1225
        "00100000", -- 0x1226
        "10010101", -- 0x1227
        "00010010", -- 0x1228
        "00100010", -- 0x1229
        "11110100", -- 0x122A
        "00010010", -- 0x122B
        "00011101", -- 0x122C
        "10100111", -- 0x122D
        "01110100", -- 0x122E
        "10000111", -- 0x122F
        "11110000", -- 0x1230
        "10010000", -- 0x1231
        "00000111", -- 0x1232
        "11001011", -- 0x1233
        "11100000", -- 0x1234
        "11111110", -- 0x1235
        "10100011", -- 0x1236
        "11100000", -- 0x1237
        "11111111", -- 0x1238
        "00010010", -- 0x1239
        "00100100", -- 0x123A
        "10010101", -- 0x123B
        "10010000", -- 0x123C
        "00010111", -- 0x123D
        "11100101", -- 0x123E
        "00010010", -- 0x123F
        "00100001", -- 0x1240
        "11001000", -- 0x1241
        "00010010", -- 0x1242
        "00100000", -- 0x1243
        "01001001", -- 0x1244
        "00100101", -- 0x1245
        "00010000", -- 0x1246
        "11111001", -- 0x1247
        "11101110", -- 0x1248
        "00110101", -- 0x1249
        "00001111", -- 0x124A
        "00010010", -- 0x124B
        "00100000", -- 0x124C
        "10010101", -- 0x124D
        "10000000", -- 0x124E
        "00010100", -- 0x124F
        "00010010", -- 0x1250
        "00100000", -- 0x1251
        "01001001", -- 0x1252
        "01111000", -- 0x1253
        "00000110", -- 0x1254
        "01111001", -- 0x1255
        "10001011", -- 0x1256
        "00101001", -- 0x1257
        "11111001", -- 0x1258
        "11101110", -- 0x1259
        "00111000", -- 0x125A
        "00010010", -- 0x125B
        "00100000", -- 0x125C
        "10010101", -- 0x125D
        "10010000", -- 0x125E
        "00000110", -- 0x125F
        "10001001", -- 0x1260
        "11100000", -- 0x1261
        "00000100", -- 0x1262
        "11110000", -- 0x1263
        "00000010", -- 0x1264
        "00100010", -- 0x1265
        "11110100", -- 0x1266
        "10001111", -- 0x1267
        "00000001", -- 0x1268
        "10001110", -- 0x1269
        "00000000", -- 0x126A
        "10010000", -- 0x126B
        "00000010", -- 0x126C
        "00001000", -- 0x126D
        "11100000", -- 0x126E
        "11111010", -- 0x126F
        "01110100", -- 0x1270
        "00100000", -- 0x1271
        "11010011", -- 0x1272
        "10011010", -- 0x1273
        "01000000", -- 0x1274
        "00100011", -- 0x1275
        "10010000", -- 0x1276
        "00000010", -- 0x1277
        "00000110", -- 0x1278
        "11100000", -- 0x1279
        "00010010", -- 0x127A
        "00011111", -- 0x127B
        "11010111", -- 0x127C
        "10001001", -- 0x127D
        "00000101", -- 0x127E
        "10001000", -- 0x127F
        "00000100", -- 0x1280
        "01111010", -- 0x1281
        "00000000", -- 0x1282
        "01111011", -- 0x1283
        "00000100", -- 0x1284
        "00010010", -- 0x1285
        "00010100", -- 0x1286
        "01111001", -- 0x1287
        "10010000", -- 0x1288
        "00000010", -- 0x1289
        "00000110", -- 0x128A
        "11100000", -- 0x128B
        "00000100", -- 0x128C
        "01010100", -- 0x128D
        "00011111", -- 0x128E
        "11110000", -- 0x128F
        "10100011", -- 0x1290
        "10100011", -- 0x1291
        "11100000", -- 0x1292
        "00000100", -- 0x1293
        "10010000", -- 0x1294
        "00000010", -- 0x1295
        "00001000", -- 0x1296
        "11110000", -- 0x1297
        "00100010", -- 0x1298
        "10001001", -- 0x1299
        "10000010", -- 0x129A
        "10001000", -- 0x129B
        "10000011", -- 0x129C
        "01111110", -- 0x129D
        "00000000", -- 0x129E
        "01111111", -- 0x129F
        "00000010", -- 0x12A0
        "00010010", -- 0x12A1
        "00100001", -- 0x12A2
        "11101011", -- 0x12A3
        "11100000", -- 0x12A4
        "00010010", -- 0x12A5
        "00100100", -- 0x12A6
        "01000010", -- 0x12A7
        "01110100", -- 0x12A8
        "00010000", -- 0x12A9
        "00010010", -- 0x12AA
        "00011111", -- 0x12AB
        "00110000", -- 0x12AC
        "00010010", -- 0x12AD
        "00100001", -- 0x12AE
        "10100100", -- 0x12AF
        "10001001", -- 0x12B0
        "00000011", -- 0x12B1
        "10001000", -- 0x12B2
        "00000010", -- 0x12B3
        "00001011", -- 0x12B4
        "10111011", -- 0x12B5
        "00000000", -- 0x12B6
        "00000001", -- 0x12B7
        "00001010", -- 0x12B8
        "10001011", -- 0x12B9
        "10000010", -- 0x12BA
        "10001010", -- 0x12BB
        "10000011", -- 0x12BC
        "11100000", -- 0x12BD
        "11111110", -- 0x12BE
        "01111111", -- 0x12BF
        "00000000", -- 0x12C0
        "00010010", -- 0x12C1
        "00100011", -- 0x12C2
        "11000000", -- 0x12C3
        "00010010", -- 0x12C4
        "00011110", -- 0x12C5
        "11110100", -- 0x12C6
        "00010010", -- 0x12C7
        "00100001", -- 0x12C8
        "10100100", -- 0x12C9
        "00010010", -- 0x12CA
        "00100100", -- 0x12CB
        "00011000", -- 0x12CC
        "00010010", -- 0x12CD
        "00011110", -- 0x12CE
        "11110100", -- 0x12CF
        "00010010", -- 0x12D0
        "00100100", -- 0x12D1
        "00010010", -- 0x12D2
        "01111111", -- 0x12D3
        "10000100", -- 0x12D4
        "00000010", -- 0x12D5
        "00010001", -- 0x12D6
        "11110101", -- 0x12D7
        "00001111", -- 0x12D8
        "10111111", -- 0x12D9
        "00000000", -- 0x12DA
        "00000001", -- 0x12DB
        "00001110", -- 0x12DC
        "10001111", -- 0x12DD
        "00001100", -- 0x12DE
        "10001110", -- 0x12DF
        "00001011", -- 0x12E0
        "10001111", -- 0x12E1
        "10000010", -- 0x12E2
        "10001110", -- 0x12E3
        "10000011", -- 0x12E4
        "11100000", -- 0x12E5
        "10110100", -- 0x12E6
        "00000001", -- 0x12E7
        "00111001", -- 0x12E8
        "10010000", -- 0x12E9
        "00000101", -- 0x12EA
        "10001001", -- 0x12EB
        "01110100", -- 0x12EC
        "01111000", -- 0x12ED
        "11110000", -- 0x12EE
        "11110000", -- 0x12EF
        "00010010", -- 0x12F0
        "00011001", -- 0x12F1
        "01001000", -- 0x12F2
        "10010000", -- 0x12F3
        "00000101", -- 0x12F4
        "10001101", -- 0x12F5
        "00010010", -- 0x12F6
        "00100001", -- 0x12F7
        "11001000", -- 0x12F8
        "00010010", -- 0x12F9
        "00100011", -- 0x12FA
        "00000110", -- 0x12FB
        "10010000", -- 0x12FC
        "00000101", -- 0x12FD
        "10010001", -- 0x12FE
        "11110000", -- 0x12FF
        "00010010", -- 0x1300
        "00100010", -- 0x1301
        "11100010", -- 0x1302
        "00010010", -- 0x1303
        "00010111", -- 0x1304
        "10001110", -- 0x1305
        "10010000", -- 0x1306
        "00000110", -- 0x1307
        "10001000", -- 0x1308
        "11110000", -- 0x1309
        "01111101", -- 0x130A
        "10000000", -- 0x130B
        "01111110", -- 0x130C
        "00000101", -- 0x130D
        "01111111", -- 0x130E
        "10010010", -- 0x130F
        "00010010", -- 0x1310
        "00011010", -- 0x1311
        "10001111", -- 0x1312
        "00010010", -- 0x1313
        "00100010", -- 0x1314
        "11100010", -- 0x1315
        "00010010", -- 0x1316
        "00011011", -- 0x1317
        "00110101", -- 0x1318
        "10010000", -- 0x1319
        "00000101", -- 0x131A
        "10001011", -- 0x131B
        "00010010", -- 0x131C
        "00011111", -- 0x131D
        "01011000", -- 0x131E
        "01110100", -- 0x131F
        "11111111", -- 0x1320
        "00100010", -- 0x1321
        "00010010", -- 0x1322
        "00100011", -- 0x1323
        "00000110", -- 0x1324
        "10110100", -- 0x1325
        "00111100", -- 0x1326
        "00000101", -- 0x1327
        "01110101", -- 0x1328
        "10000000", -- 0x1329
        "00111100", -- 0x132A
        "11100100", -- 0x132B
        "00100010", -- 0x132C
        "00010010", -- 0x132D
        "00100011", -- 0x132E
        "00000110", -- 0x132F
        "10110100", -- 0x1330
        "10111010", -- 0x1331
        "00000101", -- 0x1332
        "01110101", -- 0x1333
        "10010000", -- 0x1334
        "10111010", -- 0x1335
        "11100100", -- 0x1336
        "00100010", -- 0x1337
        "00010010", -- 0x1338
        "00100011", -- 0x1339
        "00000110", -- 0x133A
        "10110100", -- 0x133B
        "00000010", -- 0x133C
        "00000011", -- 0x133D
        "00000000", -- 0x133E
        "10000000", -- 0x133F
        "11111101", -- 0x1340
        "01110100", -- 0x1341
        "11001100", -- 0x1342
        "00100010", -- 0x1343
        "10001111", -- 0x1344
        "00011101", -- 0x1345
        "10001110", -- 0x1346
        "00011100", -- 0x1347
        "10001101", -- 0x1348
        "00011111", -- 0x1349
        "10001100", -- 0x134A
        "00011110", -- 0x134B
        "10010000", -- 0x134C
        "00000011", -- 0x134D
        "10000110", -- 0x134E
        "11100000", -- 0x134F
        "01110000", -- 0x1350
        "00011000", -- 0x1351
        "00010010", -- 0x1352
        "00011001", -- 0x1353
        "01001000", -- 0x1354
        "10010000", -- 0x1355
        "00000010", -- 0x1356
        "10001101", -- 0x1357
        "00010010", -- 0x1358
        "00100001", -- 0x1359
        "11001000", -- 0x135A
        "01111010", -- 0x135B
        "00000000", -- 0x135C
        "01111011", -- 0x135D
        "00000011", -- 0x135E
        "01111100", -- 0x135F
        "00000001", -- 0x1360
        "01111101", -- 0x1361
        "01011101", -- 0x1362
        "01111110", -- 0x1363
        "00000010", -- 0x1364
        "01111111", -- 0x1365
        "10010001", -- 0x1366
        "00010010", -- 0x1367
        "00010100", -- 0x1368
        "01111001", -- 0x1369
        "00010010", -- 0x136A
        "00100001", -- 0x136B
        "10001100", -- 0x136C
        "01111000", -- 0x136D
        "00000010", -- 0x136E
        "01111001", -- 0x136F
        "10010101", -- 0x1370
        "11101001", -- 0x1371
        "00101111", -- 0x1372
        "11111011", -- 0x1373
        "11101000", -- 0x1374
        "00111110", -- 0x1375
        "11111010", -- 0x1376
        "10001011", -- 0x1377
        "10000010", -- 0x1378
        "10001010", -- 0x1379
        "10000011", -- 0x137A
        "11100101", -- 0x137B
        "00011100", -- 0x137C
        "11110000", -- 0x137D
        "11100101", -- 0x137E
        "00011101", -- 0x137F
        "10100011", -- 0x1380
        "11110000", -- 0x1381
        "00010010", -- 0x1382
        "00100001", -- 0x1383
        "10001100", -- 0x1384
        "11101001", -- 0x1385
        "00101111", -- 0x1386
        "11111001", -- 0x1387
        "11101000", -- 0x1388
        "00111110", -- 0x1389
        "11111000", -- 0x138A
        "11101001", -- 0x138B
        "00100100", -- 0x138C
        "00000010", -- 0x138D
        "11111001", -- 0x138E
        "11100100", -- 0x138F
        "00111000", -- 0x1390
        "11111000", -- 0x1391
        "10001001", -- 0x1392
        "10000010", -- 0x1393
        "10001000", -- 0x1394
        "10000011", -- 0x1395
        "11100101", -- 0x1396
        "00011110", -- 0x1397
        "11110000", -- 0x1398
        "11100101", -- 0x1399
        "00011111", -- 0x139A
        "10100011", -- 0x139B
        "11110000", -- 0x139C
        "10010000", -- 0x139D
        "00000011", -- 0x139E
        "10000110", -- 0x139F
        "11100000", -- 0x13A0
        "00000100", -- 0x13A1
        "11110000", -- 0x13A2
        "11100000", -- 0x13A3
        "11000011", -- 0x13A4
        "10010100", -- 0x13A5
        "00111100", -- 0x13A6
        "01000000", -- 0x13A7
        "00000011", -- 0x13A8
        "00010010", -- 0x13A9
        "00010101", -- 0x13AA
        "10010000", -- 0x13AB
        "00100010", -- 0x13AC
        "10010000", -- 0x13AD
        "00000001", -- 0x13AE
        "10110101", -- 0x13AF
        "11100000", -- 0x13B0
        "10010000", -- 0x13B1
        "00000001", -- 0x13B2
        "00011110", -- 0x13B3
        "11110000", -- 0x13B4
        "10000000", -- 0x13B5
        "01010001", -- 0x13B6
        "00010010", -- 0x13B7
        "00011001", -- 0x13B8
        "01001000", -- 0x13B9
        "10010000", -- 0x13BA
        "00000001", -- 0x13BB
        "00110001", -- 0x13BC
        "00010010", -- 0x13BD
        "00100001", -- 0x13BE
        "11001000", -- 0x13BF
        "00010010", -- 0x13C0
        "00011101", -- 0x13C1
        "11111001", -- 0x13C2
        "00100100", -- 0x13C3
        "00000100", -- 0x13C4
        "00010010", -- 0x13C5
        "00100010", -- 0x13C6
        "11011001", -- 0x13C7
        "00010010", -- 0x13C8
        "00100001", -- 0x13C9
        "10111100", -- 0x13CA
        "10010000", -- 0x13CB
        "00000001", -- 0x13CC
        "00110001", -- 0x13CD
        "00010010", -- 0x13CE
        "00100011", -- 0x13CF
        "10100100", -- 0x13D0
        "01000000", -- 0x13D1
        "00110101", -- 0x13D2
        "11101001", -- 0x13D3
        "00010010", -- 0x13D4
        "00100011", -- 0x13D5
        "11011100", -- 0x13D6
        "11111010", -- 0x13D7
        "10100011", -- 0x13D8
        "11100000", -- 0x13D9
        "11111011", -- 0x13DA
        "01001010", -- 0x13DB
        "01100000", -- 0x13DC
        "00101010", -- 0x13DD
        "00010010", -- 0x13DE
        "00100100", -- 0x13DF
        "10000010", -- 0x13E0
        "11100000", -- 0x13E1
        "11111000", -- 0x13E2
        "10100011", -- 0x13E3
        "11100000", -- 0x13E4
        "11111001", -- 0x13E5
        "00010010", -- 0x13E6
        "00100100", -- 0x13E7
        "10000010", -- 0x13E8
        "00010010", -- 0x13E9
        "00100100", -- 0x13EA
        "10100010", -- 0x13EB
        "00010010", -- 0x13EC
        "00011101", -- 0x13ED
        "11111001", -- 0x13EE
        "00010010", -- 0x13EF
        "00100011", -- 0x13F0
        "11011100", -- 0x13F1
        "11111110", -- 0x13F2
        "10100011", -- 0x13F3
        "11100000", -- 0x13F4
        "11111111", -- 0x13F5
        "00010010", -- 0x13F6
        "00100100", -- 0x13F7
        "10010101", -- 0x13F8
        "10010000", -- 0x13F9
        "00000001", -- 0x13FA
        "00110001", -- 0x13FB
        "00010010", -- 0x13FC
        "00011101", -- 0x13FD
        "00010001", -- 0x13FE
        "11101001", -- 0x13FF
        "00100100", -- 0x1400
        "00000100", -- 0x1401
        "00010010", -- 0x1402
        "00100011", -- 0x1403
        "11101010", -- 0x1404
        "00010010", -- 0x1405
        "00100001", -- 0x1406
        "11001000", -- 0x1407
        "10010000", -- 0x1408
        "00000001", -- 0x1409
        "00011110", -- 0x140A
        "11100000", -- 0x140B
        "11111000", -- 0x140C
        "11100000", -- 0x140D
        "00010100", -- 0x140E
        "11110000", -- 0x140F
        "11101000", -- 0x1410
        "01110000", -- 0x1411
        "10100100", -- 0x1412
        "00100010", -- 0x1413
        "10001111", -- 0x1414
        "00000001", -- 0x1415
        "10001110", -- 0x1416
        "00000000", -- 0x1417
        "10010000", -- 0x1418
        "00000001", -- 0x1419
        "10110101", -- 0x141A
        "11100000", -- 0x141B
        "11111010", -- 0x141C
        "10000000", -- 0x141D
        "01010110", -- 0x141E
        "00011010", -- 0x141F
        "10001010", -- 0x1420
        "00000111", -- 0x1421
        "10010000", -- 0x1422
        "00000001", -- 0x1423
        "10110110", -- 0x1424
        "01110101", -- 0x1425
        "11110000", -- 0x1426
        "00001000", -- 0x1427
        "01111110", -- 0x1428
        "00000000", -- 0x1429
        "00010010", -- 0x142A
        "00011110", -- 0x142B
        "01000110", -- 0x142C
        "10000101", -- 0x142D
        "10000010", -- 0x142E
        "00010000", -- 0x142F
        "10000101", -- 0x1430
        "10000011", -- 0x1431
        "00001111", -- 0x1432
        "11100000", -- 0x1433
        "11111011", -- 0x1434
        "10100011", -- 0x1435
        "11100000", -- 0x1436
        "10110101", -- 0x1437
        "00000001", -- 0x1438
        "00111011", -- 0x1439
        "11101011", -- 0x143A
        "10110101", -- 0x143B
        "00000000", -- 0x143C
        "00110111", -- 0x143D
        "11100101", -- 0x143E
        "00010000", -- 0x143F
        "00100100", -- 0x1440
        "00000010", -- 0x1441
        "00010010", -- 0x1442
        "00100011", -- 0x1443
        "00111110", -- 0x1444
        "11101100", -- 0x1445
        "11110000", -- 0x1446
        "11101101", -- 0x1447
        "10100011", -- 0x1448
        "11110000", -- 0x1449
        "11101100", -- 0x144A
        "01001101", -- 0x144B
        "01100000", -- 0x144C
        "00001100", -- 0x144D
        "10001101", -- 0x144E
        "00000111", -- 0x144F
        "10001100", -- 0x1450
        "00000110", -- 0x1451
        "00010010", -- 0x1452
        "00000000", -- 0x1453
        "00000110", -- 0x1454
        "10010000", -- 0x1455
        "00010111", -- 0x1456
        "11011111", -- 0x1457
        "10000000", -- 0x1458
        "00001000", -- 0x1459
        "10010000", -- 0x145A
        "00010111", -- 0x145B
        "11011111", -- 0x145C
        "11100100", -- 0x145D
        "11111111", -- 0x145E
        "11111110", -- 0x145F
        "11111101", -- 0x1460
        "11111100", -- 0x1461
        "00010010", -- 0x1462
        "00100001", -- 0x1463
        "11001000", -- 0x1464
        "10010000", -- 0x1465
        "00010111", -- 0x1466
        "11011111", -- 0x1467
        "00010010", -- 0x1468
        "00100001", -- 0x1469
        "10111100", -- 0x146A
        "11100101", -- 0x146B
        "00010000", -- 0x146C
        "00100100", -- 0x146D
        "00000100", -- 0x146E
        "00010010", -- 0x146F
        "00100011", -- 0x1470
        "00111110", -- 0x1471
        "00000010", -- 0x1472
        "00100001", -- 0x1473
        "11001000", -- 0x1474
        "11101010", -- 0x1475
        "01110000", -- 0x1476
        "10100111", -- 0x1477
        "00100010", -- 0x1478
        "10010000", -- 0x1479
        "00010111", -- 0x147A
        "11100001", -- 0x147B
        "11101110", -- 0x147C
        "11110000", -- 0x147D
        "11101111", -- 0x147E
        "10100011", -- 0x147F
        "11110000", -- 0x1480
        "10010000", -- 0x1481
        "00010111", -- 0x1482
        "11100001", -- 0x1483
        "11100000", -- 0x1484
        "11111000", -- 0x1485
        "10100011", -- 0x1486
        "11100000", -- 0x1487
        "11111001", -- 0x1488
        "11101011", -- 0x1489
        "01001010", -- 0x148A
        "01100000", -- 0x148B
        "01000110", -- 0x148C
        "10101111", -- 0x148D
        "00000011", -- 0x148E
        "10010000", -- 0x148F
        "00010111", -- 0x1490
        "11100000", -- 0x1491
        "11101011", -- 0x1492
        "11110000", -- 0x1493
        "10010000", -- 0x1494
        "00010111", -- 0x1495
        "11011111", -- 0x1496
        "11101010", -- 0x1497
        "11110000", -- 0x1498
        "11101111", -- 0x1499
        "01100000", -- 0x149A
        "00001000", -- 0x149B
        "10010000", -- 0x149C
        "00010111", -- 0x149D
        "11011111", -- 0x149E
        "11100000", -- 0x149F
        "11111111", -- 0x14A0
        "00001111", -- 0x14A1
        "11101111", -- 0x14A2
        "11110000", -- 0x14A3
        "00011011", -- 0x14A4
        "10111011", -- 0x14A5
        "11111111", -- 0x14A6
        "00000001", -- 0x14A7
        "00011010", -- 0x14A8
        "10001101", -- 0x14A9
        "10000010", -- 0x14AA
        "10001100", -- 0x14AB
        "10000011", -- 0x14AC
        "11100000", -- 0x14AD
        "10001001", -- 0x14AE
        "10000010", -- 0x14AF
        "10001000", -- 0x14B0
        "10000011", -- 0x14B1
        "11110000", -- 0x14B2
        "00001001", -- 0x14B3
        "10111001", -- 0x14B4
        "00000000", -- 0x14B5
        "00000001", -- 0x14B6
        "00001000", -- 0x14B7
        "00001101", -- 0x14B8
        "10111101", -- 0x14B9
        "00000000", -- 0x14BA
        "00000001", -- 0x14BB
        "00001100", -- 0x14BC
        "10010000", -- 0x14BD
        "00010111", -- 0x14BE
        "11100000", -- 0x14BF
        "11100000", -- 0x14C0
        "11111111", -- 0x14C1
        "00011111", -- 0x14C2
        "11101111", -- 0x14C3
        "11110000", -- 0x14C4
        "10111111", -- 0x14C5
        "00000000", -- 0x14C6
        "11011100", -- 0x14C7
        "10010000", -- 0x14C8
        "00010111", -- 0x14C9
        "11011111", -- 0x14CA
        "11100000", -- 0x14CB
        "11111111", -- 0x14CC
        "00011111", -- 0x14CD
        "11101111", -- 0x14CE
        "11110000", -- 0x14CF
        "10111111", -- 0x14D0
        "00000000", -- 0x14D1
        "11010001", -- 0x14D2
        "10010000", -- 0x14D3
        "00010111", -- 0x14D4
        "11100001", -- 0x14D5
        "11100000", -- 0x14D6
        "11111110", -- 0x14D7
        "10100011", -- 0x14D8
        "11100000", -- 0x14D9
        "11111111", -- 0x14DA
        "00100010", -- 0x14DB
        "11110000", -- 0x14DC
        "10100011", -- 0x14DD
        "11100100", -- 0x14DE
        "11110000", -- 0x14DF
        "00010010", -- 0x14E0
        "00100011", -- 0x14E1
        "01111010", -- 0x14E2
        "01110100", -- 0x14E3
        "00001011", -- 0x14E4
        "11110000", -- 0x14E5
        "10100011", -- 0x14E6
        "01110100", -- 0x14E7
        "00011111", -- 0x14E8
        "11110000", -- 0x14E9
        "10100011", -- 0x14EA
        "11100100", -- 0x14EB
        "00010010", -- 0x14EC
        "00100010", -- 0x14ED
        "10111110", -- 0x14EE
        "01110100", -- 0x14EF
        "00000001", -- 0x14F0
        "11110000", -- 0x14F1
        "10100011", -- 0x14F2
        "01110100", -- 0x14F3
        "00101100", -- 0x14F4
        "00010010", -- 0x14F5
        "00100010", -- 0x14F6
        "11010000", -- 0x14F7
        "01110100", -- 0x14F8
        "00000001", -- 0x14F9
        "11110000", -- 0x14FA
        "10100011", -- 0x14FB
        "01110100", -- 0x14FC
        "11100000", -- 0x14FD
        "00010010", -- 0x14FE
        "00100011", -- 0x14FF
        "10010110", -- 0x1500
        "01110100", -- 0x1501
        "00000001", -- 0x1502
        "11110000", -- 0x1503
        "10100011", -- 0x1504
        "01110100", -- 0x1505
        "00101100", -- 0x1506
        "00010010", -- 0x1507
        "00100001", -- 0x1508
        "11010100", -- 0x1509
        "01110100", -- 0x150A
        "00010100", -- 0x150B
        "00010010", -- 0x150C
        "00100011", -- 0x150D
        "10011101", -- 0x150E
        "11100100", -- 0x150F
        "00010010", -- 0x1510
        "00100100", -- 0x1511
        "01011010", -- 0x1512
        "11100100", -- 0x1513
        "11110000", -- 0x1514
        "10100011", -- 0x1515
        "11100100", -- 0x1516
        "00010010", -- 0x1517
        "00100100", -- 0x1518
        "00000110", -- 0x1519
        "01110100", -- 0x151A
        "00001011", -- 0x151B
        "11110000", -- 0x151C
        "10100011", -- 0x151D
        "01110100", -- 0x151E
        "01110110", -- 0x151F
        "11110000", -- 0x1520
        "10100011", -- 0x1521
        "11100100", -- 0x1522
        "00010010", -- 0x1523
        "00100010", -- 0x1524
        "10111110", -- 0x1525
        "01110100", -- 0x1526
        "00000111", -- 0x1527
        "11110000", -- 0x1528
        "10100011", -- 0x1529
        "00000100", -- 0x152A
        "00010010", -- 0x152B
        "00100100", -- 0x152C
        "00000110", -- 0x152D
        "01110100", -- 0x152E
        "00001100", -- 0x152F
        "11110000", -- 0x1530
        "10100011", -- 0x1531
        "01110100", -- 0x1532
        "00110101", -- 0x1533
        "11110000", -- 0x1534
        "10100011", -- 0x1535
        "00100010", -- 0x1536
        "10111100", -- 0x1537
        "00000000", -- 0x1538
        "00000101", -- 0x1539
        "10111101", -- 0x153A
        "00000000", -- 0x153B
        "00000010", -- 0x153C
        "11010011", -- 0x153D
        "00100010", -- 0x153E
        "11000000", -- 0x153F
        "11110000", -- 0x1540
        "01110101", -- 0x1541
        "11110000", -- 0x1542
        "00000000", -- 0x1543
        "11101110", -- 0x1544
        "00110000", -- 0x1545
        "11100111", -- 0x1546
        "00001100", -- 0x1547
        "00000101", -- 0x1548
        "11110000", -- 0x1549
        "11101111", -- 0x154A
        "11110100", -- 0x154B
        "00100100", -- 0x154C
        "00000001", -- 0x154D
        "11111111", -- 0x154E
        "11101110", -- 0x154F
        "11110100", -- 0x1550
        "00110100", -- 0x1551
        "00000000", -- 0x1552
        "11111110", -- 0x1553
        "11101100", -- 0x1554
        "00110000", -- 0x1555
        "11100111", -- 0x1556
        "00010000", -- 0x1557
        "11100101", -- 0x1558
        "11110000", -- 0x1559
        "00100100", -- 0x155A
        "00000010", -- 0x155B
        "11110101", -- 0x155C
        "11110000", -- 0x155D
        "11101101", -- 0x155E
        "11110100", -- 0x155F
        "00100100", -- 0x1560
        "00000001", -- 0x1561
        "11111101", -- 0x1562
        "11101100", -- 0x1563
        "11110100", -- 0x1564
        "00110100", -- 0x1565
        "00000000", -- 0x1566
        "11111100", -- 0x1567
        "00010010", -- 0x1568
        "00001111", -- 0x1569
        "11010100", -- 0x156A
        "11100101", -- 0x156B
        "11110000", -- 0x156C
        "01100000", -- 0x156D
        "00011110", -- 0x156E
        "00110000", -- 0x156F
        "11100000", -- 0x1570
        "00001010", -- 0x1571
        "11101101", -- 0x1572
        "11110100", -- 0x1573
        "00100100", -- 0x1574
        "00000001", -- 0x1575
        "11111101", -- 0x1576
        "11101100", -- 0x1577
        "11110100", -- 0x1578
        "00110100", -- 0x1579
        "00000000", -- 0x157A
        "11111100", -- 0x157B
        "11100101", -- 0x157C
        "11110000", -- 0x157D
        "10110100", -- 0x157E
        "00000011", -- 0x157F
        "00000010", -- 0x1580
        "10000000", -- 0x1581
        "00001010", -- 0x1582
        "11101111", -- 0x1583
        "11110100", -- 0x1584
        "00100100", -- 0x1585
        "00000001", -- 0x1586
        "11111111", -- 0x1587
        "11101110", -- 0x1588
        "11110100", -- 0x1589
        "00110100", -- 0x158A
        "00000000", -- 0x158B
        "11111110", -- 0x158C
        "11010000", -- 0x158D
        "11110000", -- 0x158E
        "00100010", -- 0x158F
        "10010000", -- 0x1590
        "00000011", -- 0x1591
        "10000110", -- 0x1592
        "11100000", -- 0x1593
        "01100000", -- 0x1594
        "01010000", -- 0x1595
        "11100100", -- 0x1596
        "11111100", -- 0x1597
        "01111101", -- 0x1598
        "11111111", -- 0x1599
        "01111110", -- 0x159A
        "00000010", -- 0x159B
        "01111111", -- 0x159C
        "10001001", -- 0x159D
        "00010010", -- 0x159E
        "00010111", -- 0x159F
        "10001110", -- 0x15A0
        "10010000", -- 0x15A1
        "00000011", -- 0x15A2
        "10001000", -- 0x15A3
        "11110000", -- 0x15A4
        "01111110", -- 0x15A5
        "00000010", -- 0x15A6
        "01111111", -- 0x15A7
        "10001001", -- 0x15A8
        "00010010", -- 0x15A9
        "00011000", -- 0x15AA
        "11001111", -- 0x15AB
        "10010000", -- 0x15AC
        "00000011", -- 0x15AD
        "10000111", -- 0x15AE
        "11100000", -- 0x15AF
        "00000100", -- 0x15B0
        "11110000", -- 0x15B1
        "10010000", -- 0x15B2
        "00000011", -- 0x15B3
        "10000110", -- 0x15B4
        "11100100", -- 0x15B5
        "11110000", -- 0x15B6
        "10010000", -- 0x15B7
        "00000010", -- 0x15B8
        "10001011", -- 0x15B9
        "00010010", -- 0x15BA
        "00011111", -- 0x15BB
        "01011000", -- 0x15BC
        "01111111", -- 0x15BD
        "00000000", -- 0x15BE
        "01111000", -- 0x15BF
        "00111100", -- 0x15C0
        "10010000", -- 0x15C1
        "00000010", -- 0x15C2
        "10010101", -- 0x15C3
        "01110101", -- 0x15C4
        "11110000", -- 0x15C5
        "00000100", -- 0x15C6
        "01111110", -- 0x15C7
        "00000000", -- 0x15C8
        "00010010", -- 0x15C9
        "00011110", -- 0x15CA
        "01000110", -- 0x15CB
        "10101011", -- 0x15CC
        "10000010", -- 0x15CD
        "10101010", -- 0x15CE
        "10000011", -- 0x15CF
        "11100100", -- 0x15D0
        "11110000", -- 0x15D1
        "10100011", -- 0x15D2
        "11110000", -- 0x15D3
        "11101011", -- 0x15D4
        "00100100", -- 0x15D5
        "00000010", -- 0x15D6
        "11111011", -- 0x15D7
        "11100100", -- 0x15D8
        "00111010", -- 0x15D9
        "11111010", -- 0x15DA
        "10001011", -- 0x15DB
        "10000010", -- 0x15DC
        "10001010", -- 0x15DD
        "10000011", -- 0x15DE
        "11100100", -- 0x15DF
        "11110000", -- 0x15E0
        "10100011", -- 0x15E1
        "11110000", -- 0x15E2
        "00001111", -- 0x15E3
        "11011000", -- 0x15E4
        "11011011", -- 0x15E5
        "00100010", -- 0x15E6
        "01110101", -- 0x15E7
        "00010101", -- 0x15E8
        "00000000", -- 0x15E9
        "00010010", -- 0x15EA
        "00010110", -- 0x15EB
        "11000011", -- 0x15EC
        "00010100", -- 0x15ED
        "01100000", -- 0x15EE
        "00001000", -- 0x15EF
        "00010100", -- 0x15F0
        "01100000", -- 0x15F1
        "00010001", -- 0x15F2
        "00010100", -- 0x15F3
        "01100000", -- 0x15F4
        "00011111", -- 0x15F5
        "10000000", -- 0x15F6
        "00110010", -- 0x15F7
        "11100100", -- 0x15F8
        "11111101", -- 0x15F9
        "11111100", -- 0x15FA
        "01111110", -- 0x15FB
        "00000100", -- 0x15FC
        "01111111", -- 0x15FD
        "00010010", -- 0x15FE
        "00010010", -- 0x15FF
        "00001110", -- 0x1600
        "10011100", -- 0x1601
        "10000000", -- 0x1602
        "00100110", -- 0x1603
        "00010010", -- 0x1604
        "00100010", -- 0x1605
        "01110010", -- 0x1606
        "11111101", -- 0x1607
        "11111100", -- 0x1608
        "01111110", -- 0x1609
        "00000100", -- 0x160A
        "01111111", -- 0x160B
        "00010001", -- 0x160C
        "00010010", -- 0x160D
        "00001110", -- 0x160E
        "10011100", -- 0x160F
        "01110101", -- 0x1610
        "00010101", -- 0x1611
        "00000001", -- 0x1612
        "10000000", -- 0x1613
        "00010101", -- 0x1614
        "00010010", -- 0x1615
        "00100010", -- 0x1616
        "01110010", -- 0x1617
        "11111111", -- 0x1618
        "11111110", -- 0x1619
        "11111101", -- 0x161A
        "11111100", -- 0x161B
        "00010010", -- 0x161C
        "00100100", -- 0x161D
        "00010010", -- 0x161E
        "01111111", -- 0x161F
        "01001101", -- 0x1620
        "00010010", -- 0x1621
        "00010001", -- 0x1622
        "11110101", -- 0x1623
        "01110101", -- 0x1624
        "10011011", -- 0x1625
        "00000001", -- 0x1626
        "01110101", -- 0x1627
        "00010101", -- 0x1628
        "00000011", -- 0x1629
        "00010010", -- 0x162A
        "00011100", -- 0x162B
        "11001101", -- 0x162C
        "10010000", -- 0x162D
        "00000001", -- 0x162E
        "10100001", -- 0x162F
        "11110000", -- 0x1630
        "11100101", -- 0x1631
        "00010101", -- 0x1632
        "00100010", -- 0x1633
        "10010000", -- 0x1634
        "00010111", -- 0x1635
        "11010111", -- 0x1636
        "00010010", -- 0x1637
        "00100001", -- 0x1638
        "01110100", -- 0x1639
        "00010010", -- 0x163A
        "00011001", -- 0x163B
        "01001000", -- 0x163C
        "10010000", -- 0x163D
        "00010111", -- 0x163E
        "11010111", -- 0x163F
        "00010010", -- 0x1640
        "00011101", -- 0x1641
        "00010001", -- 0x1642
        "10010000", -- 0x1643
        "00010111", -- 0x1644
        "11011011", -- 0x1645
        "00010010", -- 0x1646
        "00100001", -- 0x1647
        "11001000", -- 0x1648
        "10000000", -- 0x1649
        "00000001", -- 0x164A
        "00000000", -- 0x164B
        "00010010", -- 0x164C
        "00100010", -- 0x164D
        "01000000", -- 0x164E
        "10010000", -- 0x164F
        "00010111", -- 0x1650
        "11011111", -- 0x1651
        "00010010", -- 0x1652
        "00100000", -- 0x1653
        "11110111", -- 0x1654
        "10010000", -- 0x1655
        "00010111", -- 0x1656
        "11100011", -- 0x1657
        "00010010", -- 0x1658
        "00100011", -- 0x1659
        "00100110", -- 0x165A
        "10010000", -- 0x165B
        "00010111", -- 0x165C
        "11100111", -- 0x165D
        "00010010", -- 0x165E
        "00100000", -- 0x165F
        "11101010", -- 0x1660
        "10010000", -- 0x1661
        "00010111", -- 0x1662
        "11011111", -- 0x1663
        "00010010", -- 0x1664
        "00011101", -- 0x1665
        "00010001", -- 0x1666
        "10010000", -- 0x1667
        "00010111", -- 0x1668
        "11100011", -- 0x1669
        "00010010", -- 0x166A
        "00011101", -- 0x166B
        "00010001", -- 0x166C
        "10010000", -- 0x166D
        "00010111", -- 0x166E
        "11100111", -- 0x166F
        "00010010", -- 0x1670
        "00011101", -- 0x1671
        "00010001", -- 0x1672
        "10010000", -- 0x1673
        "00010111", -- 0x1674
        "11011011", -- 0x1675
        "00010010", -- 0x1676
        "00100011", -- 0x1677
        "10101011", -- 0x1678
        "01000000", -- 0x1679
        "11010000", -- 0x167A
        "00100010", -- 0x167B
        "11000000", -- 0x167C
        "00000111", -- 0x167D
        "11000000", -- 0x167E
        "11100000", -- 0x167F
        "11000000", -- 0x1680
        "10000010", -- 0x1681
        "11000000", -- 0x1682
        "10000011", -- 0x1683
        "11000000", -- 0x1684
        "00000000", -- 0x1685
        "11000000", -- 0x1686
        "00000001", -- 0x1687
        "11000000", -- 0x1688
        "00000100", -- 0x1689
        "11000000", -- 0x168A
        "00000101", -- 0x168B
        "11000000", -- 0x168C
        "00000110", -- 0x168D
        "11000000", -- 0x168E
        "11010000", -- 0x168F
        "01110101", -- 0x1690
        "11010000", -- 0x1691
        "00000000", -- 0x1692
        "10010000", -- 0x1693
        "00000000", -- 0x1694
        "00000000", -- 0x1695
        "11100000", -- 0x1696
        "10010000", -- 0x1697
        "00000001", -- 0x1698
        "01100001", -- 0x1699
        "00010010", -- 0x169A
        "00100010", -- 0x169B
        "11101011", -- 0x169C
        "11100101", -- 0x169D
        "11111111", -- 0x169E
        "11110000", -- 0x169F
        "10010000", -- 0x16A0
        "00000000", -- 0x16A1
        "00000000", -- 0x16A2
        "00010010", -- 0x16A3
        "00100010", -- 0x16A4
        "01001010", -- 0x16A5
        "00010010", -- 0x16A6
        "00100011", -- 0x16A7
        "11110001", -- 0x16A8
        "10010000", -- 0x16A9
        "00000000", -- 0x16AA
        "00000000", -- 0x16AB
        "11101101", -- 0x16AC
        "11110000", -- 0x16AD
        "11010000", -- 0x16AE
        "11010000", -- 0x16AF
        "11010000", -- 0x16B0
        "00000110", -- 0x16B1
        "11010000", -- 0x16B2
        "00000101", -- 0x16B3
        "11010000", -- 0x16B4
        "00000100", -- 0x16B5
        "11010000", -- 0x16B6
        "00000001", -- 0x16B7
        "11010000", -- 0x16B8
        "00000000", -- 0x16B9
        "11010000", -- 0x16BA
        "10000011", -- 0x16BB
        "11010000", -- 0x16BC
        "10000010", -- 0x16BD
        "11010000", -- 0x16BE
        "11100000", -- 0x16BF
        "11010000", -- 0x16C0
        "00000111", -- 0x16C1
        "00110010", -- 0x16C2
        "10010000", -- 0x16C3
        "00000001", -- 0x16C4
        "00011001", -- 0x16C5
        "11100101", -- 0x16C6
        "10100000", -- 0x16C7
        "11110000", -- 0x16C8
        "11100100", -- 0x16C9
        "11111000", -- 0x16CA
        "00100000", -- 0x16CB
        "10100000", -- 0x16CC
        "00000101", -- 0x16CD
        "00100000", -- 0x16CE
        "10100010", -- 0x16CF
        "00000010", -- 0x16D0
        "01111000", -- 0x16D1
        "00000001", -- 0x16D2
        "11101000", -- 0x16D3
        "01110000", -- 0x16D4
        "00001100", -- 0x16D5
        "00100000", -- 0x16D6
        "10100000", -- 0x16D7
        "00000011", -- 0x16D8
        "00110000", -- 0x16D9
        "10100100", -- 0x16DA
        "00000110", -- 0x16DB
        "00100000", -- 0x16DC
        "10100010", -- 0x16DD
        "00000110", -- 0x16DE
        "00100000", -- 0x16DF
        "10100100", -- 0x16E0
        "00000011", -- 0x16E1
        "01110100", -- 0x16E2
        "00000001", -- 0x16E3
        "00100010", -- 0x16E4
        "11100100", -- 0x16E5
        "11111000", -- 0x16E6
        "00100000", -- 0x16E7
        "10100001", -- 0x16E8
        "00000110", -- 0x16E9
        "11100101", -- 0x16EA
        "10100000", -- 0x16EB
        "01010100", -- 0x16EC
        "00000101", -- 0x16ED
        "01100000", -- 0x16EE
        "00000110", -- 0x16EF
        "00100000", -- 0x16F0
        "10100001", -- 0x16F1
        "00000101", -- 0x16F2
        "00100000", -- 0x16F3
        "10100101", -- 0x16F4
        "00000010", -- 0x16F5
        "01111000", -- 0x16F6
        "00000001", -- 0x16F7
        "11101000", -- 0x16F8
        "01110000", -- 0x16F9
        "00000110", -- 0x16FA
        "00100000", -- 0x16FB
        "10100001", -- 0x16FC
        "00000110", -- 0x16FD
        "00100000", -- 0x16FE
        "10100101", -- 0x16FF
        "00000011", -- 0x1700
        "01110100", -- 0x1701
        "00000010", -- 0x1702
        "00100010", -- 0x1703
        "01110100", -- 0x1704
        "00000011", -- 0x1705
        "00100010", -- 0x1706
        "10001111", -- 0x1707
        "00001100", -- 0x1708
        "10001110", -- 0x1709
        "00001011", -- 0x170A
        "10010000", -- 0x170B
        "00000110", -- 0x170C
        "10001001", -- 0x170D
        "11100000", -- 0x170E
        "11111001", -- 0x170F
        "01100000", -- 0x1710
        "00110110", -- 0x1711
        "10010000", -- 0x1712
        "00000110", -- 0x1713
        "10001010", -- 0x1714
        "11100000", -- 0x1715
        "11111000", -- 0x1716
        "11101001", -- 0x1717
        "11010011", -- 0x1718
        "10011000", -- 0x1719
        "01000000", -- 0x171A
        "00001000", -- 0x171B
        "01111011", -- 0x171C
        "00100000", -- 0x171D
        "11101011", -- 0x171E
        "11000011", -- 0x171F
        "10011001", -- 0x1720
        "00101000", -- 0x1721
        "10000000", -- 0x1722
        "00000011", -- 0x1723
        "11101000", -- 0x1724
        "11000011", -- 0x1725
        "10011001", -- 0x1726
        "11111011", -- 0x1727
        "11101011", -- 0x1728
        "11111111", -- 0x1729
        "10010000", -- 0x172A
        "00000110", -- 0x172B
        "10001011", -- 0x172C
        "01110101", -- 0x172D
        "11110000", -- 0x172E
        "00001010", -- 0x172F
        "01111110", -- 0x1730
        "00000000", -- 0x1731
        "00010010", -- 0x1732
        "00011110", -- 0x1733
        "01000110", -- 0x1734
        "10101101", -- 0x1735
        "00001100", -- 0x1736
        "10101100", -- 0x1737
        "00001011", -- 0x1738
        "01111110", -- 0x1739
        "00000000", -- 0x173A
        "01111111", -- 0x173B
        "00001010", -- 0x173C
        "00010010", -- 0x173D
        "00011101", -- 0x173E
        "10000110", -- 0x173F
        "00011001", -- 0x1740
        "10010000", -- 0x1741
        "00000110", -- 0x1742
        "10001001", -- 0x1743
        "11101001", -- 0x1744
        "11110000", -- 0x1745
        "11100100", -- 0x1746
        "00100010", -- 0x1747
        "01110100", -- 0x1748
        "00000001", -- 0x1749
        "00100010", -- 0x174A
        "00010010", -- 0x174B
        "00100010", -- 0x174C
        "00000001", -- 0x174D
        "01110000", -- 0x174E
        "00111011", -- 0x174F
        "10010000", -- 0x1750
        "00011000", -- 0x1751
        "00001100", -- 0x1752
        "01110100", -- 0x1753
        "11010010", -- 0x1754
        "11110000", -- 0x1755
        "10010000", -- 0x1756
        "00000001", -- 0x1757
        "10010110", -- 0x1758
        "11100000", -- 0x1759
        "10010000", -- 0x175A
        "00011000", -- 0x175B
        "00001101", -- 0x175C
        "11110000", -- 0x175D
        "10010000", -- 0x175E
        "00000001", -- 0x175F
        "10010111", -- 0x1760
        "11100000", -- 0x1761
        "10010000", -- 0x1762
        "00011000", -- 0x1763
        "00001110", -- 0x1764
        "11110000", -- 0x1765
        "10010000", -- 0x1766
        "00000001", -- 0x1767
        "00011011", -- 0x1768
        "11100000", -- 0x1769
        "10010000", -- 0x176A
        "00011000", -- 0x176B
        "00001111", -- 0x176C
        "11110000", -- 0x176D
        "01111100", -- 0x176E
        "00000000", -- 0x176F
        "01111101", -- 0x1770
        "00000100", -- 0x1771
        "01111110", -- 0x1772
        "00011000", -- 0x1773
        "01111111", -- 0x1774
        "00001100", -- 0x1775
        "00010010", -- 0x1776
        "00010111", -- 0x1777
        "10001110", -- 0x1778
        "10010000", -- 0x1779
        "00011000", -- 0x177A
        "00010000", -- 0x177B
        "11110000", -- 0x177C
        "01111100", -- 0x177D
        "00000000", -- 0x177E
        "01111101", -- 0x177F
        "00000101", -- 0x1780
        "01111110", -- 0x1781
        "00011000", -- 0x1782
        "01111111", -- 0x1783
        "00001100", -- 0x1784
        "00010010", -- 0x1785
        "00011011", -- 0x1786
        "00110101", -- 0x1787
        "01110100", -- 0x1788
        "11111111", -- 0x1789
        "00100010", -- 0x178A
        "01110100", -- 0x178B
        "11001100", -- 0x178C
        "00100010", -- 0x178D
        "01111000", -- 0x178E
        "11111111", -- 0x178F
        "11101101", -- 0x1790
        "01001100", -- 0x1791
        "01100000", -- 0x1792
        "00111011", -- 0x1793
        "10101011", -- 0x1794
        "00000101", -- 0x1795
        "10101010", -- 0x1796
        "00000100", -- 0x1797
        "11101011", -- 0x1798
        "01100000", -- 0x1799
        "00000001", -- 0x179A
        "00001010", -- 0x179B
        "10001111", -- 0x179C
        "10000010", -- 0x179D
        "10001110", -- 0x179E
        "10000011", -- 0x179F
        "11100000", -- 0x17A0
        "11111001", -- 0x17A1
        "01101000", -- 0x17A2
        "11111000", -- 0x17A3
        "00001111", -- 0x17A4
        "10111111", -- 0x17A5
        "00000000", -- 0x17A6
        "00000001", -- 0x17A7
        "00001110", -- 0x17A8
        "11101000", -- 0x17A9
        "00000011", -- 0x17AA
        "00000011", -- 0x17AB
        "01010100", -- 0x17AC
        "11000000", -- 0x17AD
        "11111001", -- 0x17AE
        "11101000", -- 0x17AF
        "11000100", -- 0x17B0
        "01010100", -- 0x17B1
        "11110000", -- 0x17B2
        "11111100", -- 0x17B3
        "11101000", -- 0x17B4
        "11000100", -- 0x17B5
        "00000011", -- 0x17B6
        "01010100", -- 0x17B7
        "11111000", -- 0x17B8
        "01101100", -- 0x17B9
        "01101001", -- 0x17BA
        "11111001", -- 0x17BB
        "01101000", -- 0x17BC
        "11111000", -- 0x17BD
        "11000100", -- 0x17BE
        "00000011", -- 0x17BF
        "01010100", -- 0x17C0
        "00000111", -- 0x17C1
        "11111001", -- 0x17C2
        "11101000", -- 0x17C3
        "11000100", -- 0x17C4
        "01010100", -- 0x17C5
        "00001111", -- 0x17C6
        "01101001", -- 0x17C7
        "11111001", -- 0x17C8
        "01101000", -- 0x17C9
        "11111000", -- 0x17CA
        "11011011", -- 0x17CB
        "11001111", -- 0x17CC
        "11011010", -- 0x17CD
        "11001101", -- 0x17CE
        "11101000", -- 0x17CF
        "00100010", -- 0x17D0
        "10010000", -- 0x17D1
        "00000100", -- 0x17D2
        "10000100", -- 0x17D3
        "11100000", -- 0x17D4
        "01100000", -- 0x17D5
        "00111010", -- 0x17D6
        "11100100", -- 0x17D7
        "11111100", -- 0x17D8
        "01111101", -- 0x17D9
        "11111111", -- 0x17DA
        "01111110", -- 0x17DB
        "00000011", -- 0x17DC
        "01111111", -- 0x17DD
        "10001001", -- 0x17DE
        "00010010", -- 0x17DF
        "00010111", -- 0x17E0
        "10001110", -- 0x17E1
        "10010000", -- 0x17E2
        "00000100", -- 0x17E3
        "10001000", -- 0x17E4
        "11110000", -- 0x17E5
        "01111110", -- 0x17E6
        "00000011", -- 0x17E7
        "01111111", -- 0x17E8
        "10001001", -- 0x17E9
        "00010010", -- 0x17EA
        "00011000", -- 0x17EB
        "11001111", -- 0x17EC
        "10010000", -- 0x17ED
        "00000011", -- 0x17EE
        "10001011", -- 0x17EF
        "00010010", -- 0x17F0
        "00011111", -- 0x17F1
        "01011000", -- 0x17F2
        "10010000", -- 0x17F3
        "00000100", -- 0x17F4
        "10000100", -- 0x17F5
        "11100100", -- 0x17F6
        "11110000", -- 0x17F7
        "10010000", -- 0x17F8
        "00000100", -- 0x17F9
        "10000111", -- 0x17FA
        "11100000", -- 0x17FB
        "00000100", -- 0x17FC
        "11110000", -- 0x17FD
        "01111001", -- 0x17FE
        "10010100", -- 0x17FF
        "01111000", -- 0x1800
        "00000011", -- 0x1801
        "01111010", -- 0x1802
        "11110000", -- 0x1803
        "10001001", -- 0x1804
        "10000010", -- 0x1805
        "10001000", -- 0x1806
        "10000011", -- 0x1807
        "11100100", -- 0x1808
        "11110000", -- 0x1809
        "00001001", -- 0x180A
        "10111001", -- 0x180B
        "00000000", -- 0x180C
        "00000001", -- 0x180D
        "00001000", -- 0x180E
        "11011010", -- 0x180F
        "11110011", -- 0x1810
        "00100010", -- 0x1811
        "00010010", -- 0x1812
        "00100010", -- 0x1813
        "00000001", -- 0x1814
        "01100000", -- 0x1815
        "00001101", -- 0x1816
        "00010100", -- 0x1817
        "01100000", -- 0x1818
        "00101110", -- 0x1819
        "00100100", -- 0x181A
        "11111110", -- 0x181B
        "01100000", -- 0x181C
        "00010010", -- 0x181D
        "00100100", -- 0x181E
        "11111100", -- 0x181F
        "01100000", -- 0x1820
        "00011010", -- 0x1821
        "10000000", -- 0x1822
        "00101011", -- 0x1823
        "00010010", -- 0x1824
        "00100100", -- 0x1825
        "00100100", -- 0x1826
        "01100000", -- 0x1827
        "00100110", -- 0x1828
        "01111111", -- 0x1829
        "00000000", -- 0x182A
        "00010010", -- 0x182B
        "00001011", -- 0x182C
        "00110011", -- 0x182D
        "11100100", -- 0x182E
        "00100010", -- 0x182F
        "00010010", -- 0x1830
        "00100100", -- 0x1831
        "00100100", -- 0x1832
        "01100000", -- 0x1833
        "00011010", -- 0x1834
        "01111111", -- 0x1835
        "00000011", -- 0x1836
        "00010010", -- 0x1837
        "00001011", -- 0x1838
        "00110011", -- 0x1839
        "11100100", -- 0x183A
        "00100010", -- 0x183B
        "00010010", -- 0x183C
        "00100100", -- 0x183D
        "00100100", -- 0x183E
        "01100000", -- 0x183F
        "00001110", -- 0x1840
        "01111111", -- 0x1841
        "00000111", -- 0x1842
        "00010010", -- 0x1843
        "00001011", -- 0x1844
        "00110011", -- 0x1845
        "11100100", -- 0x1846
        "00100010", -- 0x1847
        "01111111", -- 0x1848
        "00000001", -- 0x1849
        "00010010", -- 0x184A
        "00001011", -- 0x184B
        "00110011", -- 0x184C
        "11100100", -- 0x184D
        "00100010", -- 0x184E
        "01110100", -- 0x184F
        "11001100", -- 0x1850
        "00100010", -- 0x1851
        "11101111", -- 0x1852
        "11110101", -- 0x1853
        "00001111", -- 0x1854
        "01100100", -- 0x1855
        "11111111", -- 0x1856
        "01100000", -- 0x1857
        "00110111", -- 0x1858
        "10010000", -- 0x1859
        "00010111", -- 0x185A
        "11010111", -- 0x185B
        "01110100", -- 0x185C
        "11001100", -- 0x185D
        "11110000", -- 0x185E
        "10100011", -- 0x185F
        "11100101", -- 0x1860
        "00001111", -- 0x1861
        "11110000", -- 0x1862
        "01111100", -- 0x1863
        "00000000", -- 0x1864
        "01111101", -- 0x1865
        "00000010", -- 0x1866
        "01111110", -- 0x1867
        "00010111", -- 0x1868
        "01111111", -- 0x1869
        "11010111", -- 0x186A
        "00010010", -- 0x186B
        "00010111", -- 0x186C
        "10001110", -- 0x186D
        "10010000", -- 0x186E
        "00010111", -- 0x186F
        "11011001", -- 0x1870
        "11110000", -- 0x1871
        "10010000", -- 0x1872
        "00010111", -- 0x1873
        "11010111", -- 0x1874
        "11100000", -- 0x1875
        "11111111", -- 0x1876
        "00010010", -- 0x1877
        "00011111", -- 0x1878
        "10110101", -- 0x1879
        "10010000", -- 0x187A
        "00010111", -- 0x187B
        "11011000", -- 0x187C
        "11100000", -- 0x187D
        "11111111", -- 0x187E
        "00010010", -- 0x187F
        "00011111", -- 0x1880
        "10110101", -- 0x1881
        "10010000", -- 0x1882
        "00010111", -- 0x1883
        "11011001", -- 0x1884
        "11100000", -- 0x1885
        "11111111", -- 0x1886
        "00010010", -- 0x1887
        "00011111", -- 0x1888
        "10110101", -- 0x1889
        "10010000", -- 0x188A
        "00000000", -- 0x188B
        "00000011", -- 0x188C
        "11100101", -- 0x188D
        "00001111", -- 0x188E
        "11110000", -- 0x188F
        "00100010", -- 0x1890
        "10010000", -- 0x1891
        "00000010", -- 0x1892
        "00001000", -- 0x1893
        "11100000", -- 0x1894
        "11111000", -- 0x1895
        "10010000", -- 0x1896
        "00000010", -- 0x1897
        "00000110", -- 0x1898
        "11100000", -- 0x1899
        "11111011", -- 0x189A
        "01111010", -- 0x189B
        "00000000", -- 0x189C
        "11000011", -- 0x189D
        "10011000", -- 0x189E
        "11111101", -- 0x189F
        "11100100", -- 0x18A0
        "10011010", -- 0x18A1
        "00110000", -- 0x18A2
        "11100111", -- 0x18A3
        "00001100", -- 0x18A4
        "11101000", -- 0x18A5
        "11000011", -- 0x18A6
        "10011011", -- 0x18A7
        "11111011", -- 0x18A8
        "01111101", -- 0x18A9
        "00100000", -- 0x18AA
        "11101101", -- 0x18AB
        "11000011", -- 0x18AC
        "10011011", -- 0x18AD
        "11111011", -- 0x18AE
        "10000000", -- 0x18AF
        "00000010", -- 0x18B0
        "10001101", -- 0x18B1
        "00000011", -- 0x18B2
        "11101000", -- 0x18B3
        "01100000", -- 0x18B4
        "00011000", -- 0x18B5
        "11101011", -- 0x18B6
        "00010010", -- 0x18B7
        "00011111", -- 0x18B8
        "11010111", -- 0x18B9
        "00010010", -- 0x18BA
        "00001101", -- 0x18BB
        "01010011", -- 0x18BC
        "10010000", -- 0x18BD
        "00000010", -- 0x18BE
        "00001000", -- 0x18BF
        "11100000", -- 0x18C0
        "00010100", -- 0x18C1
        "11110000", -- 0x18C2
        "11100000", -- 0x18C3
        "11010011", -- 0x18C4
        "10010100", -- 0x18C5
        "00100000", -- 0x18C6
        "01000000", -- 0x18C7
        "00000101", -- 0x18C8
        "10010000", -- 0x18C9
        "00000010", -- 0x18CA
        "00001000", -- 0x18CB
        "11100100", -- 0x18CC
        "11110000", -- 0x18CD
        "00100010", -- 0x18CE
        "10001111", -- 0x18CF
        "00000101", -- 0x18D0
        "10001110", -- 0x18D1
        "00000100", -- 0x18D2
        "10010000", -- 0x18D3
        "00000111", -- 0x18D4
        "11001111", -- 0x18D5
        "11100000", -- 0x18D6
        "11111000", -- 0x18D7
        "01110100", -- 0x18D8
        "00010000", -- 0x18D9
        "11010011", -- 0x18DA
        "10011000", -- 0x18DB
        "01000000", -- 0x18DC
        "00011110", -- 0x18DD
        "10010000", -- 0x18DE
        "00000111", -- 0x18DF
        "11001101", -- 0x18E0
        "00010010", -- 0x18E1
        "00100001", -- 0x18E2
        "00000100", -- 0x18E3
        "01111010", -- 0x18E4
        "00000001", -- 0x18E5
        "01111011", -- 0x18E6
        "00000000", -- 0x18E7
        "00010010", -- 0x18E8
        "00010100", -- 0x18E9
        "01111001", -- 0x18EA
        "10010000", -- 0x18EB
        "00000111", -- 0x18EC
        "11001101", -- 0x18ED
        "11100000", -- 0x18EE
        "00000100", -- 0x18EF
        "01010100", -- 0x18F0
        "00001111", -- 0x18F1
        "11110000", -- 0x18F2
        "10100011", -- 0x18F3
        "10100011", -- 0x18F4
        "11100000", -- 0x18F5
        "00000100", -- 0x18F6
        "10010000", -- 0x18F7
        "00000111", -- 0x18F8
        "11001111", -- 0x18F9
        "11110000", -- 0x18FA
        "00100010", -- 0x18FB
        "11100100", -- 0x18FC
        "11111111", -- 0x18FD
        "11111110", -- 0x18FE
        "11111101", -- 0x18FF
        "11111100", -- 0x1900
        "10010000", -- 0x1901
        "00010111", -- 0x1902
        "11101001", -- 0x1903
        "00010010", -- 0x1904
        "00100001", -- 0x1905
        "11001000", -- 0x1906
        "01111111", -- 0x1907
        "10000000", -- 0x1908
        "00000010", -- 0x1909
        "00010001", -- 0x190A
        "11110101", -- 0x190B
        "10010000", -- 0x190C
        "00000111", -- 0x190D
        "11001111", -- 0x190E
        "11100000", -- 0x190F
        "11111100", -- 0x1910
        "10010000", -- 0x1911
        "00000111", -- 0x1912
        "11001101", -- 0x1913
        "11100000", -- 0x1914
        "11111001", -- 0x1915
        "01111000", -- 0x1916
        "00000000", -- 0x1917
        "11000011", -- 0x1918
        "10011100", -- 0x1919
        "11111011", -- 0x191A
        "11100100", -- 0x191B
        "10011000", -- 0x191C
        "00110000", -- 0x191D
        "11100111", -- 0x191E
        "00001001", -- 0x191F
        "01111011", -- 0x1920
        "00010000", -- 0x1921
        "11101011", -- 0x1922
        "11000011", -- 0x1923
        "10011100", -- 0x1924
        "00101001", -- 0x1925
        "11111001", -- 0x1926
        "10000000", -- 0x1927
        "00000010", -- 0x1928
        "10001011", -- 0x1929
        "00000001", -- 0x192A
        "11101001", -- 0x192B
        "11111000", -- 0x192C
        "11101100", -- 0x192D
        "01100000", -- 0x192E
        "00010111", -- 0x192F
        "01111001", -- 0x1930
        "00000000", -- 0x1931
        "11101001", -- 0x1932
        "00100100", -- 0x1933
        "11010000", -- 0x1934
        "11111101", -- 0x1935
        "11101000", -- 0x1936
        "00110100", -- 0x1937
        "00000111", -- 0x1938
        "11111100", -- 0x1939
        "01111010", -- 0x193A
        "00000001", -- 0x193B
        "01111011", -- 0x193C
        "00000000", -- 0x193D
        "00010010", -- 0x193E
        "00010100", -- 0x193F
        "01111001", -- 0x1940
        "10010000", -- 0x1941
        "00000111", -- 0x1942
        "11001111", -- 0x1943
        "11100000", -- 0x1944
        "00010100", -- 0x1945
        "11110000", -- 0x1946
        "00100010", -- 0x1947
        "01110101", -- 0x1948
        "11001100", -- 0x1949
        "00000001", -- 0x194A
        "00010010", -- 0x194B
        "00100010", -- 0x194C
        "01000000", -- 0x194D
        "10010000", -- 0x194E
        "00010111", -- 0x194F
        "11110001", -- 0x1950
        "00010010", -- 0x1951
        "00100000", -- 0x1952
        "11110111", -- 0x1953
        "10010000", -- 0x1954
        "00010111", -- 0x1955
        "11110101", -- 0x1956
        "00010010", -- 0x1957
        "00100011", -- 0x1958
        "00100110", -- 0x1959
        "10010000", -- 0x195A
        "00010111", -- 0x195B
        "11111001", -- 0x195C
        "00010010", -- 0x195D
        "00100000", -- 0x195E
        "11101010", -- 0x195F
        "10010000", -- 0x1960
        "00010111", -- 0x1961
        "11110001", -- 0x1962
        "00010010", -- 0x1963
        "00011101", -- 0x1964
        "00010001", -- 0x1965
        "10010000", -- 0x1966
        "00010111", -- 0x1967
        "11110101", -- 0x1968
        "00010010", -- 0x1969
        "00011101", -- 0x196A
        "00010001", -- 0x196B
        "10010000", -- 0x196C
        "00010111", -- 0x196D
        "11111001", -- 0x196E
        "00010010", -- 0x196F
        "00011101", -- 0x1970
        "00010001", -- 0x1971
        "10010000", -- 0x1972
        "00010111", -- 0x1973
        "11101101", -- 0x1974
        "00010010", -- 0x1975
        "00100001", -- 0x1976
        "11001000", -- 0x1977
        "01110101", -- 0x1978
        "11001100", -- 0x1979
        "00000000", -- 0x197A
        "10010000", -- 0x197B
        "00010111", -- 0x197C
        "11101101", -- 0x197D
        "00000010", -- 0x197E
        "00100001", -- 0x197F
        "10111100", -- 0x1980
        "10001111", -- 0x1981
        "00010001", -- 0x1982
        "10010000", -- 0x1983
        "00000100", -- 0x1984
        "10000100", -- 0x1985
        "11100000", -- 0x1986
        "01110000", -- 0x1987
        "00010100", -- 0x1988
        "00010010", -- 0x1989
        "00011001", -- 0x198A
        "01001000", -- 0x198B
        "10010000", -- 0x198C
        "00000011", -- 0x198D
        "10001101", -- 0x198E
        "00010010", -- 0x198F
        "00100001", -- 0x1990
        "11001000", -- 0x1991
        "00010010", -- 0x1992
        "00100000", -- 0x1993
        "11011101", -- 0x1994
        "11101000", -- 0x1995
        "00100101", -- 0x1996
        "11100000", -- 0x1997
        "01001001", -- 0x1998
        "10010000", -- 0x1999
        "00000011", -- 0x199A
        "10010001", -- 0x199B
        "11110000", -- 0x199C
        "10010000", -- 0x199D
        "00000100", -- 0x199E
        "10000100", -- 0x199F
        "11100000", -- 0x19A0
        "10010000", -- 0x19A1
        "00000011", -- 0x19A2
        "10010100", -- 0x19A3
        "00010010", -- 0x19A4
        "00100010", -- 0x19A5
        "11101011", -- 0x19A6
        "11100101", -- 0x19A7
        "00010001", -- 0x19A8
        "11110000", -- 0x19A9
        "10010000", -- 0x19AA
        "00000100", -- 0x19AB
        "10000100", -- 0x19AC
        "11100000", -- 0x19AD
        "00000100", -- 0x19AE
        "11110000", -- 0x19AF
        "11100000", -- 0x19B0
        "11000011", -- 0x19B1
        "10010100", -- 0x19B2
        "11110000", -- 0x19B3
        "01000000", -- 0x19B4
        "00000011", -- 0x19B5
        "00010010", -- 0x19B6
        "00010111", -- 0x19B7
        "11010001", -- 0x19B8
        "00100010", -- 0x19B9
        "00000001", -- 0x19BA
        "00000011", -- 0x19BB
        "00010001", -- 0x19BC
        "00000010", -- 0x19BD
        "00000010", -- 0x19BE
        "10101010", -- 0x19BF
        "00000100", -- 0x19C0
        "00000010", -- 0x19C1
        "11001111", -- 0x19C2
        "00000101", -- 0x19C3
        "00000010", -- 0x19C4
        "11010111", -- 0x19C5
        "00000110", -- 0x19C6
        "00000010", -- 0x19C7
        "00101100", -- 0x19C8
        "00000111", -- 0x19C9
        "00000010", -- 0x19CA
        "00011000", -- 0x19CB
        "00001000", -- 0x19CC
        "00000001", -- 0x19CD
        "11110001", -- 0x19CE
        "00001001", -- 0x19CF
        "00000010", -- 0x19D0
        "00110111", -- 0x19D1
        "00001010", -- 0x19D2
        "00000010", -- 0x19D3
        "11100110", -- 0x19D4
        "00001011", -- 0x19D5
        "00000010", -- 0x19D6
        "01111000", -- 0x19D7
        "00001100", -- 0x19D8
        "00000010", -- 0x19D9
        "01010001", -- 0x19DA
        "00001101", -- 0x19DB
        "00000010", -- 0x19DC
        "10010111", -- 0x19DD
        "00001110", -- 0x19DE
        "00000010", -- 0x19DF
        "11111100", -- 0x19E0
        "00001111", -- 0x19E1
        "00000010", -- 0x19E2
        "11101100", -- 0x19E3
        "00010000", -- 0x19E4
        "00000001", -- 0x19E5
        "11111010", -- 0x19E6
        "00010001", -- 0x19E7
        "00000001", -- 0x19E8
        "10010100", -- 0x19E9
        "10100000", -- 0x19EA
        "00000001", -- 0x19EB
        "11000100", -- 0x19EC
        "10100001", -- 0x19ED
        "00000001", -- 0x19EE
        "11011110", -- 0x19EF
        "10100010", -- 0x19F0
        "00000010", -- 0x19F1
        "00000100", -- 0x19F2
        "01110101", -- 0x19F3
        "11100101", -- 0x19F4
        "00000000", -- 0x19F5
        "01010011", -- 0x19F6
        "11101101", -- 0x19F7
        "00111111", -- 0x19F8
        "01000011", -- 0x19F9
        "11101101", -- 0x19FA
        "10000000", -- 0x19FB
        "01010011", -- 0x19FC
        "11101101", -- 0x19FD
        "11001111", -- 0x19FE
        "01000011", -- 0x19FF
        "11101101", -- 0x1A00
        "00100000", -- 0x1A01
        "01110101", -- 0x1A02
        "10110000", -- 0x1A03
        "00000000", -- 0x1A04
        "01010011", -- 0x1A05
        "11010101", -- 0x1A06
        "11001111", -- 0x1A07
        "01000011", -- 0x1A08
        "11010101", -- 0x1A09
        "00100000", -- 0x1A0A
        "01010011", -- 0x1A0B
        "11010101", -- 0x1A0C
        "11110011", -- 0x1A0D
        "01000011", -- 0x1A0E
        "11010101", -- 0x1A0F
        "00001000", -- 0x1A10
        "01110101", -- 0x1A11
        "11010100", -- 0x1A12
        "00000000", -- 0x1A13
        "01110101", -- 0x1A14
        "11111101", -- 0x1A15
        "00100110", -- 0x1A16
        "01110101", -- 0x1A17
        "11110101", -- 0x1A18
        "00100101", -- 0x1A19
        "00010010", -- 0x1A1A
        "00010101", -- 0x1A1B
        "11100111", -- 0x1A1C
        "11100100", -- 0x1A1D
        "01111111", -- 0x1A1E
        "10000000", -- 0x1A1F
        "01111110", -- 0x1A20
        "00100101", -- 0x1A21
        "11111101", -- 0x1A22
        "11111100", -- 0x1A23
        "00010010", -- 0x1A24
        "00001101", -- 0x1A25
        "11111001", -- 0x1A26
        "01110101", -- 0x1A27
        "10100000", -- 0x1A28
        "00000010", -- 0x1A29
        "00100010", -- 0x1A2A
        "10010000", -- 0x1A2B
        "00000100", -- 0x1A2C
        "10000100", -- 0x1A2D
        "11100000", -- 0x1A2E
        "10110100", -- 0x1A2F
        "00000001", -- 0x1A30
        "00011011", -- 0x1A31
        "00010010", -- 0x1A32
        "00011001", -- 0x1A33
        "01001000", -- 0x1A34
        "10010000", -- 0x1A35
        "00000000", -- 0x1A36
        "00001100", -- 0x1A37
        "00010010", -- 0x1A38
        "00011010", -- 0x1A39
        "11100100", -- 0x1A3A
        "10010000", -- 0x1A3B
        "00011000", -- 0x1A3C
        "00100101", -- 0x1A3D
        "00010010", -- 0x1A3E
        "00100001", -- 0x1A3F
        "11001000", -- 0x1A40
        "10010000", -- 0x1A41
        "00011000", -- 0x1A42
        "00100111", -- 0x1A43
        "00010010", -- 0x1A44
        "00100100", -- 0x1A45
        "01110011", -- 0x1A46
        "10010000", -- 0x1A47
        "00000011", -- 0x1A48
        "10010010", -- 0x1A49
        "00010010", -- 0x1A4A
        "00100100", -- 0x1A4B
        "01010100", -- 0x1A4C
        "10010000", -- 0x1A4D
        "00000001", -- 0x1A4E
        "10010110", -- 0x1A4F
        "11100000", -- 0x1A50
        "11111111", -- 0x1A51
        "00010010", -- 0x1A52
        "00011001", -- 0x1A53
        "10000001", -- 0x1A54
        "00010010", -- 0x1A55
        "00011001", -- 0x1A56
        "01001000", -- 0x1A57
        "10010000", -- 0x1A58
        "00000000", -- 0x1A59
        "00001100", -- 0x1A5A
        "00000010", -- 0x1A5B
        "00100001", -- 0x1A5C
        "11001000", -- 0x1A5D
        "11000000", -- 0x1A5E
        "10000011", -- 0x1A5F
        "11000000", -- 0x1A60
        "10000010", -- 0x1A61
        "11100000", -- 0x1A62
        "11000000", -- 0x1A63
        "11100000", -- 0x1A64
        "10100011", -- 0x1A65
        "11100000", -- 0x1A66
        "11000000", -- 0x1A67
        "11100000", -- 0x1A68
        "10100011", -- 0x1A69
        "11100000", -- 0x1A6A
        "11000000", -- 0x1A6B
        "11100000", -- 0x1A6C
        "10100011", -- 0x1A6D
        "11100000", -- 0x1A6E
        "11000000", -- 0x1A6F
        "11100000", -- 0x1A70
        "00010010", -- 0x1A71
        "00010000", -- 0x1A72
        "01101011", -- 0x1A73
        "11010000", -- 0x1A74
        "11100000", -- 0x1A75
        "11111111", -- 0x1A76
        "11010000", -- 0x1A77
        "11100000", -- 0x1A78
        "11111110", -- 0x1A79
        "11010000", -- 0x1A7A
        "11100000", -- 0x1A7B
        "11111101", -- 0x1A7C
        "11010000", -- 0x1A7D
        "11100000", -- 0x1A7E
        "11111100", -- 0x1A7F
        "11010000", -- 0x1A80
        "10000010", -- 0x1A81
        "11010000", -- 0x1A82
        "10000011", -- 0x1A83
        "11110000", -- 0x1A84
        "10100011", -- 0x1A85
        "11101101", -- 0x1A86
        "11110000", -- 0x1A87
        "10100011", -- 0x1A88
        "11101110", -- 0x1A89
        "11110000", -- 0x1A8A
        "10100011", -- 0x1A8B
        "11101111", -- 0x1A8C
        "11110000", -- 0x1A8D
        "00100010", -- 0x1A8E
        "10001111", -- 0x1A8F
        "00001110", -- 0x1A90
        "10001110", -- 0x1A91
        "00001101", -- 0x1A92
        "10001101", -- 0x1A93
        "00000001", -- 0x1A94
        "01110101", -- 0x1A95
        "11110000", -- 0x1A96
        "00000000", -- 0x1A97
        "11101001", -- 0x1A98
        "01100000", -- 0x1A99
        "00011111", -- 0x1A9A
        "11110101", -- 0x1A9B
        "00001111", -- 0x1A9C
        "00011001", -- 0x1A9D
        "10101111", -- 0x1A9E
        "11110000", -- 0x1A9F
        "00010010", -- 0x1AA0
        "00011100", -- 0x1AA1
        "00011100", -- 0x1AA2
        "10000101", -- 0x1AA3
        "00001110", -- 0x1AA4
        "10000010", -- 0x1AA5
        "10000101", -- 0x1AA6
        "00001101", -- 0x1AA7
        "10000011", -- 0x1AA8
        "11110000", -- 0x1AA9
        "00000101", -- 0x1AAA
        "00001110", -- 0x1AAB
        "11100101", -- 0x1AAC
        "00001110", -- 0x1AAD
        "01110000", -- 0x1AAE
        "00000010", -- 0x1AAF
        "00000101", -- 0x1AB0
        "00001101", -- 0x1AB1
        "00000101", -- 0x1AB2
        "11110000", -- 0x1AB3
        "00010101", -- 0x1AB4
        "00001111", -- 0x1AB5
        "11100101", -- 0x1AB6
        "00001111", -- 0x1AB7
        "01110000", -- 0x1AB8
        "11100011", -- 0x1AB9
        "00100010", -- 0x1ABA
        "00010010", -- 0x1ABB
        "00100010", -- 0x1ABC
        "00000001", -- 0x1ABD
        "01110000", -- 0x1ABE
        "00011011", -- 0x1ABF
        "10010000", -- 0x1AC0
        "00000111", -- 0x1AC1
        "11001111", -- 0x1AC2
        "11100000", -- 0x1AC3
        "01100000", -- 0x1AC4
        "00011011", -- 0x1AC5
        "01111110", -- 0x1AC6
        "00000100", -- 0x1AC7
        "01111111", -- 0x1AC8
        "10001001", -- 0x1AC9
        "00010010", -- 0x1ACA
        "00011001", -- 0x1ACB
        "00001100", -- 0x1ACC
        "01111100", -- 0x1ACD
        "00000001", -- 0x1ACE
        "01111101", -- 0x1ACF
        "00000000", -- 0x1AD0
        "01111110", -- 0x1AD1
        "00000100", -- 0x1AD2
        "01111111", -- 0x1AD3
        "10001001", -- 0x1AD4
        "00010010", -- 0x1AD5
        "00011011", -- 0x1AD6
        "00110101", -- 0x1AD7
        "01110100", -- 0x1AD8
        "11111111", -- 0x1AD9
        "00100010", -- 0x1ADA
        "10010000", -- 0x1ADB
        "00000100", -- 0x1ADC
        "10001001", -- 0x1ADD
        "11100000", -- 0x1ADE
        "01110000", -- 0x1ADF
        "11101100", -- 0x1AE0
        "01110100", -- 0x1AE1
        "11001100", -- 0x1AE2
        "00100010", -- 0x1AE3
        "11000000", -- 0x1AE4
        "00000000", -- 0x1AE5
        "11000000", -- 0x1AE6
        "00000001", -- 0x1AE7
        "11000000", -- 0x1AE8
        "00000010", -- 0x1AE9
        "11000000", -- 0x1AEA
        "00000011", -- 0x1AEB
        "11100000", -- 0x1AEC
        "11111000", -- 0x1AED
        "10100011", -- 0x1AEE
        "11100000", -- 0x1AEF
        "11111001", -- 0x1AF0
        "10100011", -- 0x1AF1
        "11100000", -- 0x1AF2
        "11111010", -- 0x1AF3
        "10100011", -- 0x1AF4
        "11100000", -- 0x1AF5
        "11111011", -- 0x1AF6
        "11000011", -- 0x1AF7
        "11101111", -- 0x1AF8
        "10011011", -- 0x1AF9
        "11111111", -- 0x1AFA
        "11101110", -- 0x1AFB
        "10011010", -- 0x1AFC
        "11111110", -- 0x1AFD
        "11101101", -- 0x1AFE
        "10011001", -- 0x1AFF
        "11111101", -- 0x1B00
        "11101100", -- 0x1B01
        "10011000", -- 0x1B02
        "11111100", -- 0x1B03
        "11010000", -- 0x1B04
        "00000011", -- 0x1B05
        "11010000", -- 0x1B06
        "00000010", -- 0x1B07
        "11010000", -- 0x1B08
        "00000001", -- 0x1B09
        "11010000", -- 0x1B0A
        "00000000", -- 0x1B0B
        "00100010", -- 0x1B0C
        "10010000", -- 0x1B0D
        "00000001", -- 0x1B0E
        "00111101", -- 0x1B0F
        "11100100", -- 0x1B10
        "11110000", -- 0x1B11
        "10010000", -- 0x1B12
        "00000001", -- 0x1B13
        "01000101", -- 0x1B14
        "11100100", -- 0x1B15
        "11110000", -- 0x1B16
        "10010000", -- 0x1B17
        "00000001", -- 0x1B18
        "00111110", -- 0x1B19
        "11100100", -- 0x1B1A
        "11110000", -- 0x1B1B
        "01110100", -- 0x1B1C
        "00001010", -- 0x1B1D
        "10100011", -- 0x1B1E
        "11110000", -- 0x1B1F
        "10100011", -- 0x1B20
        "11100100", -- 0x1B21
        "11110000", -- 0x1B22
        "10100011", -- 0x1B23
        "11110000", -- 0x1B24
        "10010000", -- 0x1B25
        "00000001", -- 0x1B26
        "01000010", -- 0x1B27
        "11100100", -- 0x1B28
        "11110000", -- 0x1B29
        "10100011", -- 0x1B2A
        "01110100", -- 0x1B2B
        "11101111", -- 0x1B2C
        "11110000", -- 0x1B2D
        "10100011", -- 0x1B2E
        "01110100", -- 0x1B2F
        "00000001", -- 0x1B30
        "11110000", -- 0x1B31
        "00000010", -- 0x1B32
        "00100010", -- 0x1B33
        "01010100", -- 0x1B34
        "10001111", -- 0x1B35
        "00000001", -- 0x1B36
        "10001110", -- 0x1B37
        "00000000", -- 0x1B38
        "11101101", -- 0x1B39
        "01001100", -- 0x1B3A
        "01100000", -- 0x1B3B
        "00011111", -- 0x1B3C
        "10101011", -- 0x1B3D
        "00000101", -- 0x1B3E
        "10101010", -- 0x1B3F
        "00000100", -- 0x1B40
        "11101011", -- 0x1B41
        "01100000", -- 0x1B42
        "00000001", -- 0x1B43
        "00001010", -- 0x1B44
        "00011101", -- 0x1B45
        "10111101", -- 0x1B46
        "11111111", -- 0x1B47
        "00000001", -- 0x1B48
        "00011100", -- 0x1B49
        "10001001", -- 0x1B4A
        "10000010", -- 0x1B4B
        "10001000", -- 0x1B4C
        "10000011", -- 0x1B4D
        "11100000", -- 0x1B4E
        "11111111", -- 0x1B4F
        "00010010", -- 0x1B50
        "00011111", -- 0x1B51
        "10110101", -- 0x1B52
        "00001001", -- 0x1B53
        "10111001", -- 0x1B54
        "00000000", -- 0x1B55
        "00000001", -- 0x1B56
        "00001000", -- 0x1B57
        "11011011", -- 0x1B58
        "11101011", -- 0x1B59
        "11011010", -- 0x1B5A
        "11101001", -- 0x1B5B
        "00100010", -- 0x1B5C
        "11000011", -- 0x1B5D
        "11000000", -- 0x1B5E
        "10000011", -- 0x1B5F
        "11000000", -- 0x1B60
        "10000010", -- 0x1B61
        "11100000", -- 0x1B62
        "11000000", -- 0x1B63
        "11100000", -- 0x1B64
        "10100011", -- 0x1B65
        "11100000", -- 0x1B66
        "11000000", -- 0x1B67
        "11100000", -- 0x1B68
        "10100011", -- 0x1B69
        "11100000", -- 0x1B6A
        "11000000", -- 0x1B6B
        "11100000", -- 0x1B6C
        "10100011", -- 0x1B6D
        "11100000", -- 0x1B6E
        "11000000", -- 0x1B6F
        "11100000", -- 0x1B70
        "00010010", -- 0x1B71
        "00011110", -- 0x1B72
        "10100001", -- 0x1B73
        "11010000", -- 0x1B74
        "10000010", -- 0x1B75
        "11010000", -- 0x1B76
        "10000011", -- 0x1B77
        "11101100", -- 0x1B78
        "11110000", -- 0x1B79
        "10100011", -- 0x1B7A
        "11101101", -- 0x1B7B
        "11110000", -- 0x1B7C
        "10100011", -- 0x1B7D
        "11101110", -- 0x1B7E
        "11110000", -- 0x1B7F
        "10100011", -- 0x1B80
        "11101111", -- 0x1B81
        "11110000", -- 0x1B82
        "00100010", -- 0x1B83
        "11000000", -- 0x1B84
        "10000011", -- 0x1B85
        "11000000", -- 0x1B86
        "10000010", -- 0x1B87
        "11100000", -- 0x1B88
        "11111101", -- 0x1B89
        "10100011", -- 0x1B8A
        "11100000", -- 0x1B8B
        "11111110", -- 0x1B8C
        "10100011", -- 0x1B8D
        "11100000", -- 0x1B8E
        "11111111", -- 0x1B8F
        "10100011", -- 0x1B90
        "11100000", -- 0x1B91
        "00100100", -- 0x1B92
        "11111111", -- 0x1B93
        "11110000", -- 0x1B94
        "11001111", -- 0x1B95
        "00110100", -- 0x1B96
        "11111111", -- 0x1B97
        "11001110", -- 0x1B98
        "00110100", -- 0x1B99
        "11111111", -- 0x1B9A
        "11001101", -- 0x1B9B
        "00110100", -- 0x1B9C
        "11111111", -- 0x1B9D
        "11111100", -- 0x1B9E
        "11010000", -- 0x1B9F
        "10000010", -- 0x1BA0
        "11010000", -- 0x1BA1
        "10000011", -- 0x1BA2
        "11110000", -- 0x1BA3
        "11101101", -- 0x1BA4
        "10100011", -- 0x1BA5
        "11110000", -- 0x1BA6
        "11101110", -- 0x1BA7
        "10100011", -- 0x1BA8
        "11110000", -- 0x1BA9
        "00100010", -- 0x1BAA
        "10001111", -- 0x1BAB
        "00001100", -- 0x1BAC
        "10001110", -- 0x1BAD
        "00001011", -- 0x1BAE
        "10001101", -- 0x1BAF
        "00000001", -- 0x1BB0
        "01111010", -- 0x1BB1
        "00000000", -- 0x1BB2
        "11101001", -- 0x1BB3
        "01100000", -- 0x1BB4
        "00011010", -- 0x1BB5
        "11111011", -- 0x1BB6
        "00011001", -- 0x1BB7
        "10000101", -- 0x1BB8
        "00001100", -- 0x1BB9
        "10000010", -- 0x1BBA
        "10000101", -- 0x1BBB
        "00001011", -- 0x1BBC
        "10000011", -- 0x1BBD
        "11100000", -- 0x1BBE
        "11111101", -- 0x1BBF
        "10001010", -- 0x1BC0
        "00000111", -- 0x1BC1
        "00010010", -- 0x1BC2
        "00011111", -- 0x1BC3
        "01111111", -- 0x1BC4
        "00000101", -- 0x1BC5
        "00001100", -- 0x1BC6
        "11100101", -- 0x1BC7
        "00001100", -- 0x1BC8
        "01110000", -- 0x1BC9
        "00000010", -- 0x1BCA
        "00000101", -- 0x1BCB
        "00001011", -- 0x1BCC
        "00001010", -- 0x1BCD
        "11011011", -- 0x1BCE
        "11100111", -- 0x1BCF
        "00100010", -- 0x1BD0
        "11000000", -- 0x1BD1
        "10000011", -- 0x1BD2
        "11000000", -- 0x1BD3
        "10000010", -- 0x1BD4
        "11100000", -- 0x1BD5
        "11000000", -- 0x1BD6
        "11100000", -- 0x1BD7
        "10100011", -- 0x1BD8
        "11100000", -- 0x1BD9
        "11000000", -- 0x1BDA
        "11100000", -- 0x1BDB
        "10100011", -- 0x1BDC
        "11100000", -- 0x1BDD
        "11000000", -- 0x1BDE
        "11100000", -- 0x1BDF
        "10100011", -- 0x1BE0
        "11100000", -- 0x1BE1
        "11000000", -- 0x1BE2
        "11100000", -- 0x1BE3
        "00010010", -- 0x1BE4
        "00011111", -- 0x1BE5
        "00001000", -- 0x1BE6
        "11010000", -- 0x1BE7
        "10000010", -- 0x1BE8
        "11010000", -- 0x1BE9
        "10000011", -- 0x1BEA
        "11101100", -- 0x1BEB
        "11110000", -- 0x1BEC
        "10100011", -- 0x1BED
        "11101101", -- 0x1BEE
        "11110000", -- 0x1BEF
        "10100011", -- 0x1BF0
        "11101110", -- 0x1BF1
        "11110000", -- 0x1BF2
        "10100011", -- 0x1BF3
        "11101111", -- 0x1BF4
        "11110000", -- 0x1BF5
        "00100010", -- 0x1BF6
        "11001010", -- 0x1BF7
        "11000000", -- 0x1BF8
        "11100000", -- 0x1BF9
        "11100100", -- 0x1BFA
        "10010011", -- 0x1BFB
        "01101010", -- 0x1BFC
        "10100011", -- 0x1BFD
        "01100000", -- 0x1BFE
        "00001001", -- 0x1BFF
        "10100011", -- 0x1C00
        "10100011", -- 0x1C01
        "11010101", -- 0x1C02
        "11110000", -- 0x1C03
        "11110101", -- 0x1C04
        "11010000", -- 0x1C05
        "11100000", -- 0x1C06
        "11111010", -- 0x1C07
        "00100010", -- 0x1C08
        "11100100", -- 0x1C09
        "10010011", -- 0x1C0A
        "11111010", -- 0x1C0B
        "10100011", -- 0x1C0C
        "11100100", -- 0x1C0D
        "10010011", -- 0x1C0E
        "11110101", -- 0x1C0F
        "10000010", -- 0x1C10
        "10001010", -- 0x1C11
        "10000011", -- 0x1C12
        "11010000", -- 0x1C13
        "11100000", -- 0x1C14
        "11111010", -- 0x1C15
        "11010000", -- 0x1C16
        "11100000", -- 0x1C17
        "11010000", -- 0x1C18
        "11100000", -- 0x1C19
        "11100100", -- 0x1C1A
        "01110011", -- 0x1C1B
        "10101000", -- 0x1C1C
        "11101110", -- 0x1C1D
        "10001111", -- 0x1C1E
        "11111110", -- 0x1C1F
        "01110101", -- 0x1C20
        "11101110", -- 0x1C21
        "00000000", -- 0x1C22
        "01111000", -- 0x1C23
        "00000000", -- 0x1C24
        "10000000", -- 0x1C25
        "00000001", -- 0x1C26
        "00000000", -- 0x1C27
        "11100101", -- 0x1C28
        "11101110", -- 0x1C29
        "01010100", -- 0x1C2A
        "00000001", -- 0x1C2B
        "11111011", -- 0x1C2C
        "11100100", -- 0x1C2D
        "11111010", -- 0x1C2E
        "01001011", -- 0x1C2F
        "01110000", -- 0x1C30
        "11110101", -- 0x1C31
        "10101000", -- 0x1C32
        "11101110", -- 0x1C33
        "11100100", -- 0x1C34
        "11111110", -- 0x1C35
        "11111101", -- 0x1C36
        "11111100", -- 0x1C37
        "01111111", -- 0x1C38
        "00000001", -- 0x1C39
        "00010010", -- 0x1C3A
        "00010110", -- 0x1C3B
        "00110100", -- 0x1C3C
        "11100101", -- 0x1C3D
        "11110110", -- 0x1C3E
        "00100010", -- 0x1C3F
        "11000000", -- 0x1C40
        "11100000", -- 0x1C41
        "11100101", -- 0x1C42
        "10000001", -- 0x1C43
        "00010100", -- 0x1C44
        "00010100", -- 0x1C45
        "00010100", -- 0x1C46
        "11001000", -- 0x1C47
        "11000110", -- 0x1C48
        "00011000", -- 0x1C49
        "11001001", -- 0x1C4A
        "11000110", -- 0x1C4B
        "00011000", -- 0x1C4C
        "11001001", -- 0x1C4D
        "11000110", -- 0x1C4E
        "00011000", -- 0x1C4F
        "11001001", -- 0x1C50
        "11000110", -- 0x1C51
        "00011000", -- 0x1C52
        "11001001", -- 0x1C53
        "11000110", -- 0x1C54
        "00011000", -- 0x1C55
        "11001001", -- 0x1C56
        "11000110", -- 0x1C57
        "00001000", -- 0x1C58
        "00001000", -- 0x1C59
        "00001000", -- 0x1C5A
        "00001000", -- 0x1C5B
        "11000110", -- 0x1C5C
        "00001000", -- 0x1C5D
        "11001001", -- 0x1C5E
        "11000110", -- 0x1C5F
        "11001000", -- 0x1C60
        "11010000", -- 0x1C61
        "11100000", -- 0x1C62
        "00100010", -- 0x1C63
        "11000000", -- 0x1C64
        "11100000", -- 0x1C65
        "11100101", -- 0x1C66
        "10000001", -- 0x1C67
        "00010100", -- 0x1C68
        "00010100", -- 0x1C69
        "00010100", -- 0x1C6A
        "11001000", -- 0x1C6B
        "11000110", -- 0x1C6C
        "00011000", -- 0x1C6D
        "11001001", -- 0x1C6E
        "11000110", -- 0x1C6F
        "00011000", -- 0x1C70
        "00011000", -- 0x1C71
        "00011000", -- 0x1C72
        "00011000", -- 0x1C73
        "11000110", -- 0x1C74
        "00001000", -- 0x1C75
        "11001001", -- 0x1C76
        "11000110", -- 0x1C77
        "00001000", -- 0x1C78
        "11001001", -- 0x1C79
        "11000110", -- 0x1C7A
        "00001000", -- 0x1C7B
        "11001001", -- 0x1C7C
        "11000110", -- 0x1C7D
        "00001000", -- 0x1C7E
        "11001001", -- 0x1C7F
        "11000110", -- 0x1C80
        "00001000", -- 0x1C81
        "11001001", -- 0x1C82
        "11000110", -- 0x1C83
        "11001000", -- 0x1C84
        "11010000", -- 0x1C85
        "11100000", -- 0x1C86
        "00100010", -- 0x1C87
        "11000000", -- 0x1C88
        "00000000", -- 0x1C89
        "11000000", -- 0x1C8A
        "00000001", -- 0x1C8B
        "11000000", -- 0x1C8C
        "00000010", -- 0x1C8D
        "11100000", -- 0x1C8E
        "11111000", -- 0x1C8F
        "10100011", -- 0x1C90
        "11100000", -- 0x1C91
        "11111001", -- 0x1C92
        "10100011", -- 0x1C93
        "11100000", -- 0x1C94
        "11111010", -- 0x1C95
        "10100011", -- 0x1C96
        "11100000", -- 0x1C97
        "11000011", -- 0x1C98
        "10011111", -- 0x1C99
        "11111111", -- 0x1C9A
        "11101010", -- 0x1C9B
        "10011110", -- 0x1C9C
        "11111110", -- 0x1C9D
        "11101001", -- 0x1C9E
        "10011101", -- 0x1C9F
        "11111101", -- 0x1CA0
        "11101000", -- 0x1CA1
        "10011100", -- 0x1CA2
        "11111100", -- 0x1CA3
        "11010000", -- 0x1CA4
        "00000010", -- 0x1CA5
        "11010000", -- 0x1CA6
        "00000001", -- 0x1CA7
        "11010000", -- 0x1CA8
        "00000000", -- 0x1CA9
        "00100010", -- 0x1CAA
        "11100101", -- 0x1CAB
        "00001100", -- 0x1CAC
        "00100100", -- 0x1CAD
        "00000010", -- 0x1CAE
        "00010010", -- 0x1CAF
        "00100000", -- 0x1CB0
        "11000001", -- 0x1CB1
        "00010010", -- 0x1CB2
        "00100001", -- 0x1CB3
        "11001000", -- 0x1CB4
        "00010010", -- 0x1CB5
        "00100100", -- 0x1CB6
        "00011000", -- 0x1CB7
        "01110100", -- 0x1CB8
        "00001000", -- 0x1CB9
        "00010010", -- 0x1CBA
        "00011111", -- 0x1CBB
        "00110000", -- 0x1CBC
        "10010000", -- 0x1CBD
        "00010111", -- 0x1CBE
        "11010011", -- 0x1CBF
        "00010010", -- 0x1CC0
        "00100001", -- 0x1CC1
        "11001000", -- 0x1CC2
        "11100101", -- 0x1CC3
        "00001100", -- 0x1CC4
        "00100100", -- 0x1CC5
        "00000011", -- 0x1CC6
        "00010010", -- 0x1CC7
        "00100000", -- 0x1CC8
        "11000001", -- 0x1CC9
        "00000010", -- 0x1CCA
        "00011011", -- 0x1CCB
        "11010001", -- 0x1CCC
        "01111101", -- 0x1CCD
        "00001011", -- 0x1CCE
        "01111110", -- 0x1CCF
        "00011000", -- 0x1CD0
        "01111111", -- 0x1CD1
        "00010001", -- 0x1CD2
        "00010010", -- 0x1CD3
        "00011010", -- 0x1CD4
        "10001111", -- 0x1CD5
        "01111100", -- 0x1CD6
        "00000000", -- 0x1CD7
        "01111101", -- 0x1CD8
        "00001010", -- 0x1CD9
        "01111110", -- 0x1CDA
        "00011000", -- 0x1CDB
        "01111111", -- 0x1CDC
        "00010001", -- 0x1CDD
        "00010010", -- 0x1CDE
        "00010111", -- 0x1CDF
        "10001110", -- 0x1CE0
        "11111000", -- 0x1CE1
        "10010000", -- 0x1CE2
        "00011000", -- 0x1CE3
        "00011011", -- 0x1CE4
        "11100000", -- 0x1CE5
        "10110101", -- 0x1CE6
        "00000000", -- 0x1CE7
        "00000011", -- 0x1CE8
        "01110100", -- 0x1CE9
        "01011010", -- 0x1CEA
        "00100010", -- 0x1CEB
        "01110100", -- 0x1CEC
        "10100101", -- 0x1CED
        "00100010", -- 0x1CEE
        "11110000", -- 0x1CEF
        "10010000", -- 0x1CF0
        "00000001", -- 0x1CF1
        "01011000", -- 0x1CF2
        "11100100", -- 0x1CF3
        "11110000", -- 0x1CF4
        "10100011", -- 0x1CF5
        "11110000", -- 0x1CF6
        "10101101", -- 0x1CF7
        "00001110", -- 0x1CF8
        "10101100", -- 0x1CF9
        "00001101", -- 0x1CFA
        "01111010", -- 0x1CFB
        "00000000", -- 0x1CFC
        "01111011", -- 0x1CFD
        "00000011", -- 0x1CFE
        "01111110", -- 0x1CFF
        "00000001", -- 0x1D00
        "01111111", -- 0x1D01
        "01011101", -- 0x1D02
        "00010010", -- 0x1D03
        "00010100", -- 0x1D04
        "01111001", -- 0x1D05
        "01111100", -- 0x1D06
        "00000000", -- 0x1D07
        "01111101", -- 0x1D08
        "01100100", -- 0x1D09
        "01111110", -- 0x1D0A
        "00000100", -- 0x1D0B
        "01111111", -- 0x1D0C
        "11001101", -- 0x1D0D
        "00000010", -- 0x1D0E
        "00010100", -- 0x1D0F
        "00010100", -- 0x1D10
        "11000000", -- 0x1D11
        "00000000", -- 0x1D12
        "11000000", -- 0x1D13
        "00000001", -- 0x1D14
        "11000000", -- 0x1D15
        "00000010", -- 0x1D16
        "11100000", -- 0x1D17
        "11111000", -- 0x1D18
        "10100011", -- 0x1D19
        "11100000", -- 0x1D1A
        "11111001", -- 0x1D1B
        "10100011", -- 0x1D1C
        "11100000", -- 0x1D1D
        "11111010", -- 0x1D1E
        "10100011", -- 0x1D1F
        "11100000", -- 0x1D20
        "00101111", -- 0x1D21
        "11111111", -- 0x1D22
        "11101010", -- 0x1D23
        "00111110", -- 0x1D24
        "11111110", -- 0x1D25
        "11101001", -- 0x1D26
        "00111101", -- 0x1D27
        "11111101", -- 0x1D28
        "11101000", -- 0x1D29
        "00111100", -- 0x1D2A
        "11111100", -- 0x1D2B
        "11010000", -- 0x1D2C
        "00000010", -- 0x1D2D
        "11010000", -- 0x1D2E
        "00000001", -- 0x1D2F
        "11010000", -- 0x1D30
        "00000000", -- 0x1D31
        "00100010", -- 0x1D32
        "10010000", -- 0x1D33
        "00000001", -- 0x1D34
        "10000101", -- 0x1D35
        "01110100", -- 0x1D36
        "01010101", -- 0x1D37
        "11110000", -- 0x1D38
        "10100011", -- 0x1D39
        "01110100", -- 0x1D3A
        "00110100", -- 0x1D3B
        "11110000", -- 0x1D3C
        "10010000", -- 0x1D3D
        "00000001", -- 0x1D3E
        "10110011", -- 0x1D3F
        "01110100", -- 0x1D40
        "00011101", -- 0x1D41
        "11110000", -- 0x1D42
        "10010000", -- 0x1D43
        "00000001", -- 0x1D44
        "10000111", -- 0x1D45
        "11100100", -- 0x1D46
        "11110000", -- 0x1D47
        "10100011", -- 0x1D48
        "11110000", -- 0x1D49
        "10010000", -- 0x1D4A
        "00000001", -- 0x1D4B
        "10110010", -- 0x1D4C
        "01110100", -- 0x1D4D
        "00000001", -- 0x1D4E
        "11110000", -- 0x1D4F
        "00100010", -- 0x1D50
        "10010000", -- 0x1D51
        "00000000", -- 0x1D52
        "00000010", -- 0x1D53
        "00010010", -- 0x1D54
        "00100010", -- 0x1D55
        "01001010", -- 0x1D56
        "00010010", -- 0x1D57
        "00100000", -- 0x1D58
        "10000110", -- 0x1D59
        "10010000", -- 0x1D5A
        "00011000", -- 0x1D5B
        "00100001", -- 0x1D5C
        "11110000", -- 0x1D5D
        "00010010", -- 0x1D5E
        "00100011", -- 0x1D5F
        "10110010", -- 0x1D60
        "00100100", -- 0x1D61
        "00000010", -- 0x1D62
        "11111111", -- 0x1D63
        "11100100", -- 0x1D64
        "00111000", -- 0x1D65
        "11111110", -- 0x1D66
        "00010010", -- 0x1D67
        "00100000", -- 0x1D68
        "10000110", -- 0x1D69
        "10010000", -- 0x1D6A
        "00011000", -- 0x1D6B
        "00100010", -- 0x1D6C
        "11110000", -- 0x1D6D
        "00100010", -- 0x1D6E
        "11100000", -- 0x1D6F
        "10100011", -- 0x1D70
        "11001100", -- 0x1D71
        "11000101", -- 0x1D72
        "10000011", -- 0x1D73
        "11001101", -- 0x1D74
        "11000101", -- 0x1D75
        "10000010", -- 0x1D76
        "11001100", -- 0x1D77
        "11110000", -- 0x1D78
        "10100011", -- 0x1D79
        "11001101", -- 0x1D7A
        "11000101", -- 0x1D7B
        "10000011", -- 0x1D7C
        "11001100", -- 0x1D7D
        "11000101", -- 0x1D7E
        "10000010", -- 0x1D7F
        "11001101", -- 0x1D80
        "11101111", -- 0x1D81
        "01110000", -- 0x1D82
        "00000001", -- 0x1D83
        "00011110", -- 0x1D84
        "00011111", -- 0x1D85
        "11101110", -- 0x1D86
        "01001111", -- 0x1D87
        "01110000", -- 0x1D88
        "11100101", -- 0x1D89
        "00100010", -- 0x1D8A
        "00010010", -- 0x1D8B
        "00100010", -- 0x1D8C
        "10101100", -- 0x1D8D
        "01110101", -- 0x1D8E
        "10110000", -- 0x1D8F
        "00000000", -- 0x1D90
        "10000101", -- 0x1D91
        "00001110", -- 0x1D92
        "10000010", -- 0x1D93
        "10000101", -- 0x1D94
        "00001101", -- 0x1D95
        "10000011", -- 0x1D96
        "11100000", -- 0x1D97
        "10010000", -- 0x1D98
        "00000001", -- 0x1D99
        "01010001", -- 0x1D9A
        "11110000", -- 0x1D9B
        "11100101", -- 0x1D9C
        "00001100", -- 0x1D9D
        "00100100", -- 0x1D9E
        "00000010", -- 0x1D9F
        "11111001", -- 0x1DA0
        "11100100", -- 0x1DA1
        "00110101", -- 0x1DA2
        "00001011", -- 0x1DA3
        "00000010", -- 0x1DA4
        "00100100", -- 0x1DA5
        "10011001", -- 0x1DA6
        "00010010", -- 0x1DA7
        "00011001", -- 0x1DA8
        "01001000", -- 0x1DA9
        "10010000", -- 0x1DAA
        "00010111", -- 0x1DAB
        "11100001", -- 0x1DAC
        "00010010", -- 0x1DAD
        "00100001", -- 0x1DAE
        "11001000", -- 0x1DAF
        "10010000", -- 0x1DB0
        "00000001", -- 0x1DB1
        "00011101", -- 0x1DB2
        "11100000", -- 0x1DB3
        "11111000", -- 0x1DB4
        "10010000", -- 0x1DB5
        "00010111", -- 0x1DB6
        "11011111", -- 0x1DB7
        "11110000", -- 0x1DB8
        "00001000", -- 0x1DB9
        "10010000", -- 0x1DBA
        "00000001", -- 0x1DBB
        "00011101", -- 0x1DBC
        "11101000", -- 0x1DBD
        "11110000", -- 0x1DBE
        "10010000", -- 0x1DBF
        "00010111", -- 0x1DC0
        "11100000", -- 0x1DC1
        "00100010", -- 0x1DC2
        "11100000", -- 0x1DC3
        "11000000", -- 0x1DC4
        "11100000", -- 0x1DC5
        "10100011", -- 0x1DC6
        "11100000", -- 0x1DC7
        "11000000", -- 0x1DC8
        "11100000", -- 0x1DC9
        "10100011", -- 0x1DCA
        "11100000", -- 0x1DCB
        "11000000", -- 0x1DCC
        "11100000", -- 0x1DCD
        "10100011", -- 0x1DCE
        "11100000", -- 0x1DCF
        "11000000", -- 0x1DD0
        "11100000", -- 0x1DD1
        "00010010", -- 0x1DD2
        "00010000", -- 0x1DD3
        "01101011", -- 0x1DD4
        "11010000", -- 0x1DD5
        "00000111", -- 0x1DD6
        "11010000", -- 0x1DD7
        "00000110", -- 0x1DD8
        "11010000", -- 0x1DD9
        "00000101", -- 0x1DDA
        "11010000", -- 0x1DDB
        "00000100", -- 0x1DDC
        "00100010", -- 0x1DDD
        "11100000", -- 0x1DDE
        "11000000", -- 0x1DDF
        "11100000", -- 0x1DE0
        "10100011", -- 0x1DE1
        "11100000", -- 0x1DE2
        "11000000", -- 0x1DE3
        "11100000", -- 0x1DE4
        "10100011", -- 0x1DE5
        "11100000", -- 0x1DE6
        "11000000", -- 0x1DE7
        "11100000", -- 0x1DE8
        "10100011", -- 0x1DE9
        "11100000", -- 0x1DEA
        "11000000", -- 0x1DEB
        "11100000", -- 0x1DEC
        "00010010", -- 0x1DED
        "00010000", -- 0x1DEE
        "01101011", -- 0x1DEF
        "11010000", -- 0x1DF0
        "11100000", -- 0x1DF1
        "11010000", -- 0x1DF2
        "11100000", -- 0x1DF3
        "11010000", -- 0x1DF4
        "11100000", -- 0x1DF5
        "11010000", -- 0x1DF6
        "11100000", -- 0x1DF7
        "00100010", -- 0x1DF8
        "10010000", -- 0x1DF9
        "00000001", -- 0x1DFA
        "10110110", -- 0x1DFB
        "10101001", -- 0x1DFC
        "10000010", -- 0x1DFD
        "10101000", -- 0x1DFE
        "10000011", -- 0x1DFF
        "10010000", -- 0x1E00
        "00000001", -- 0x1E01
        "00011110", -- 0x1E02
        "11100000", -- 0x1E03
        "00010010", -- 0x1E04
        "00100100", -- 0x1E05
        "10000010", -- 0x1E06
        "01110101", -- 0x1E07
        "11110000", -- 0x1E08
        "00001000", -- 0x1E09
        "00010010", -- 0x1E0A
        "00100001", -- 0x1E0B
        "01011100", -- 0x1E0C
        "10101001", -- 0x1E0D
        "10000010", -- 0x1E0E
        "10101000", -- 0x1E0F
        "10000011", -- 0x1E10
        "11101001", -- 0x1E11
        "00100010", -- 0x1E12
        "11000000", -- 0x1E13
        "11100000", -- 0x1E14
        "11000000", -- 0x1E15
        "10000010", -- 0x1E16
        "11000000", -- 0x1E17
        "10000011", -- 0x1E18
        "11000000", -- 0x1E19
        "11010000", -- 0x1E1A
        "01110101", -- 0x1E1B
        "11010000", -- 0x1E1C
        "00000000", -- 0x1E1D
        "10010000", -- 0x1E1E
        "00000000", -- 0x1E1F
        "00000001", -- 0x1E20
        "01110100", -- 0x1E21
        "00000001", -- 0x1E22
        "11110000", -- 0x1E23
        "11010000", -- 0x1E24
        "11010000", -- 0x1E25
        "11010000", -- 0x1E26
        "10000011", -- 0x1E27
        "11010000", -- 0x1E28
        "10000010", -- 0x1E29
        "11010000", -- 0x1E2A
        "11100000", -- 0x1E2B
        "00110010", -- 0x1E2C
        "00100100", -- 0x1E2D
        "11111111", -- 0x1E2E
        "10110011", -- 0x1E2F
        "11100100", -- 0x1E30
        "00110011", -- 0x1E31
        "11111111", -- 0x1E32
        "01111101", -- 0x1E33
        "00000100", -- 0x1E34
        "01111110", -- 0x1E35
        "00000000", -- 0x1E36
        "00010010", -- 0x1E37
        "00100000", -- 0x1E38
        "00001001", -- 0x1E39
        "11101111", -- 0x1E3A
        "00100100", -- 0x1E3B
        "00010000", -- 0x1E3C
        "01000010", -- 0x1E3D
        "11101101", -- 0x1E3E
        "01010011", -- 0x1E3F
        "11101101", -- 0x1E40
        "00111111", -- 0x1E41
        "01000011", -- 0x1E42
        "11101101", -- 0x1E43
        "01000000", -- 0x1E44
        "00100010", -- 0x1E45
        "11000000", -- 0x1E46
        "11110000", -- 0x1E47
        "11101111", -- 0x1E48
        "10100100", -- 0x1E49
        "00100101", -- 0x1E4A
        "10000010", -- 0x1E4B
        "11110101", -- 0x1E4C
        "10000010", -- 0x1E4D
        "11100101", -- 0x1E4E
        "10000011", -- 0x1E4F
        "00110101", -- 0x1E50
        "11110000", -- 0x1E51
        "11110101", -- 0x1E52
        "10000011", -- 0x1E53
        "11010000", -- 0x1E54
        "11110000", -- 0x1E55
        "11101110", -- 0x1E56
        "10100100", -- 0x1E57
        "00100101", -- 0x1E58
        "10000011", -- 0x1E59
        "11110101", -- 0x1E5A
        "10000011", -- 0x1E5B
        "00100010", -- 0x1E5C
        "10010000", -- 0x1E5D
        "00000010", -- 0x1E5E
        "10001010", -- 0x1E5F
        "01110100", -- 0x1E60
        "01010101", -- 0x1E61
        "11110000", -- 0x1E62
        "10010000", -- 0x1E63
        "00000010", -- 0x1E64
        "10001001", -- 0x1E65
        "00010010", -- 0x1E66
        "00100010", -- 0x1E67
        "10010000", -- 0x1E68
        "10010000", -- 0x1E69
        "00000011", -- 0x1E6A
        "10000111", -- 0x1E6B
        "11100100", -- 0x1E6C
        "11110000", -- 0x1E6D
        "10010000", -- 0x1E6E
        "00000011", -- 0x1E6F
        "10000110", -- 0x1E70
        "11100100", -- 0x1E71
        "11110000", -- 0x1E72
        "00100010", -- 0x1E73
        "10010000", -- 0x1E74
        "00000011", -- 0x1E75
        "10001010", -- 0x1E76
        "01110100", -- 0x1E77
        "11001100", -- 0x1E78
        "11110000", -- 0x1E79
        "10010000", -- 0x1E7A
        "00000011", -- 0x1E7B
        "10001001", -- 0x1E7C
        "00010010", -- 0x1E7D
        "00100010", -- 0x1E7E
        "10010000", -- 0x1E7F
        "10010000", -- 0x1E80
        "00000100", -- 0x1E81
        "10000111", -- 0x1E82
        "11100100", -- 0x1E83
        "11110000", -- 0x1E84
        "10010000", -- 0x1E85
        "00000100", -- 0x1E86
        "10000100", -- 0x1E87
        "11100100", -- 0x1E88
        "11110000", -- 0x1E89
        "00100010", -- 0x1E8A
        "11100000", -- 0x1E8B
        "11001110", -- 0x1E8C
        "10100011", -- 0x1E8D
        "11100000", -- 0x1E8E
        "11001111", -- 0x1E8F
        "11111101", -- 0x1E90
        "00010010", -- 0x1E91
        "00100000", -- 0x1E92
        "00001001", -- 0x1E93
        "11101111", -- 0x1E94
        "11110000", -- 0x1E95
        "11100101", -- 0x1E96
        "10000010", -- 0x1E97
        "01110000", -- 0x1E98
        "00000010", -- 0x1E99
        "00010101", -- 0x1E9A
        "10000011", -- 0x1E9B
        "00010101", -- 0x1E9C
        "10000010", -- 0x1E9D
        "11101110", -- 0x1E9E
        "11110000", -- 0x1E9F
        "00100010", -- 0x1EA0
        "00010010", -- 0x1EA1
        "00011100", -- 0x1EA2
        "01100100", -- 0x1EA3
        "11010000", -- 0x1EA4
        "11100000", -- 0x1EA5
        "11000011", -- 0x1EA6
        "10011111", -- 0x1EA7
        "11111111", -- 0x1EA8
        "11010000", -- 0x1EA9
        "11100000", -- 0x1EAA
        "10011110", -- 0x1EAB
        "11111110", -- 0x1EAC
        "11010000", -- 0x1EAD
        "11100000", -- 0x1EAE
        "10011101", -- 0x1EAF
        "11111101", -- 0x1EB0
        "11010000", -- 0x1EB1
        "11100000", -- 0x1EB2
        "10011100", -- 0x1EB3
        "11111100", -- 0x1EB4
        "00100010", -- 0x1EB5
        "11000000", -- 0x1EB6
        "11110000", -- 0x1EB7
        "11101101", -- 0x1EB8
        "10001111", -- 0x1EB9
        "11110000", -- 0x1EBA
        "10100100", -- 0x1EBB
        "11001111", -- 0x1EBC
        "11000101", -- 0x1EBD
        "11110000", -- 0x1EBE
        "11001100", -- 0x1EBF
        "10100100", -- 0x1EC0
        "00101100", -- 0x1EC1
        "11001110", -- 0x1EC2
        "10001101", -- 0x1EC3
        "11110000", -- 0x1EC4
        "10100100", -- 0x1EC5
        "00101110", -- 0x1EC6
        "11111110", -- 0x1EC7
        "11010000", -- 0x1EC8
        "11110000", -- 0x1EC9
        "00100010", -- 0x1ECA
        "00010010", -- 0x1ECB
        "00100011", -- 0x1ECC
        "11010101", -- 0x1ECD
        "10010000", -- 0x1ECE
        "00000001", -- 0x1ECF
        "01011100", -- 0x1ED0
        "11100000", -- 0x1ED1
        "00000100", -- 0x1ED2
        "11110000", -- 0x1ED3
        "11100000", -- 0x1ED4
        "00010010", -- 0x1ED5
        "00100100", -- 0x1ED6
        "01000010", -- 0x1ED7
        "00010010", -- 0x1ED8
        "00100100", -- 0x1ED9
        "00010010", -- 0x1EDA
        "01111111", -- 0x1EDB
        "00001110", -- 0x1EDC
        "00000010", -- 0x1EDD
        "00010001", -- 0x1EDE
        "11110101", -- 0x1EDF
        "00010010", -- 0x1EE0
        "00011001", -- 0x1EE1
        "11110011", -- 0x1EE2
        "00010010", -- 0x1EE3
        "00100100", -- 0x1EE4
        "00111100", -- 0x1EE5
        "10010000", -- 0x1EE6
        "00000001", -- 0x1EE7
        "01001110", -- 0x1EE8
        "00010010", -- 0x1EE9
        "00011111", -- 0x1EEA
        "01011000", -- 0x1EEB
        "00010010", -- 0x1EEC
        "00100011", -- 0x1EED
        "01010110", -- 0x1EEE
        "01111111", -- 0x1EEF
        "00000001", -- 0x1EF0
        "00000010", -- 0x1EF1
        "00010001", -- 0x1EF2
        "11110101", -- 0x1EF3
        "00010010", -- 0x1EF4
        "00011100", -- 0x1EF5
        "01100100", -- 0x1EF6
        "11010000", -- 0x1EF7
        "11100000", -- 0x1EF8
        "01001111", -- 0x1EF9
        "11111111", -- 0x1EFA
        "11010000", -- 0x1EFB
        "11100000", -- 0x1EFC
        "01001110", -- 0x1EFD
        "11111110", -- 0x1EFE
        "11010000", -- 0x1EFF
        "11100000", -- 0x1F00
        "01001101", -- 0x1F01
        "11111101", -- 0x1F02
        "11010000", -- 0x1F03
        "11100000", -- 0x1F04
        "01001100", -- 0x1F05
        "11111100", -- 0x1F06
        "00100010", -- 0x1F07
        "00010010", -- 0x1F08
        "00011100", -- 0x1F09
        "01100100", -- 0x1F0A
        "11010000", -- 0x1F0B
        "11100000", -- 0x1F0C
        "00101111", -- 0x1F0D
        "11111111", -- 0x1F0E
        "11010000", -- 0x1F0F
        "11100000", -- 0x1F10
        "00111110", -- 0x1F11
        "11111110", -- 0x1F12
        "11010000", -- 0x1F13
        "11100000", -- 0x1F14
        "00111101", -- 0x1F15
        "11111101", -- 0x1F16
        "11010000", -- 0x1F17
        "11100000", -- 0x1F18
        "00111100", -- 0x1F19
        "11111100", -- 0x1F1A
        "00100010", -- 0x1F1B
        "01010100", -- 0x1F1C
        "00011111", -- 0x1F1D
        "01100000", -- 0x1F1E
        "00001111", -- 0x1F1F
        "11001100", -- 0x1F20
        "11000011", -- 0x1F21
        "00010011", -- 0x1F22
        "11001101", -- 0x1F23
        "00010011", -- 0x1F24
        "11001101", -- 0x1F25
        "11001110", -- 0x1F26
        "00010011", -- 0x1F27
        "11001110", -- 0x1F28
        "11001111", -- 0x1F29
        "00010011", -- 0x1F2A
        "11001111", -- 0x1F2B
        "11011100", -- 0x1F2C
        "11110011", -- 0x1F2D
        "11111100", -- 0x1F2E
        "00100010", -- 0x1F2F
        "01010100", -- 0x1F30
        "00011111", -- 0x1F31
        "01100000", -- 0x1F32
        "00001111", -- 0x1F33
        "11001111", -- 0x1F34
        "00100101", -- 0x1F35
        "11100000", -- 0x1F36
        "11001110", -- 0x1F37
        "00110011", -- 0x1F38
        "11001110", -- 0x1F39
        "11001101", -- 0x1F3A
        "00110011", -- 0x1F3B
        "11001101", -- 0x1F3C
        "11001100", -- 0x1F3D
        "00110011", -- 0x1F3E
        "11001100", -- 0x1F3F
        "11011111", -- 0x1F40
        "11110011", -- 0x1F41
        "11111111", -- 0x1F42
        "00100010", -- 0x1F43
        "01111111", -- 0x1F44
        "00001000", -- 0x1F45
        "00010010", -- 0x1F46
        "00011110", -- 0x1F47
        "10001011", -- 0x1F48
        "11100101", -- 0x1F49
        "00001100", -- 0x1F4A
        "00100100", -- 0x1F4B
        "00000011", -- 0x1F4C
        "11111001", -- 0x1F4D
        "11100100", -- 0x1F4E
        "00110101", -- 0x1F4F
        "00001011", -- 0x1F50
        "00010010", -- 0x1F51
        "00100100", -- 0x1F52
        "10011001", -- 0x1F53
        "11111111", -- 0x1F54
        "01111110", -- 0x1F55
        "00000000", -- 0x1F56
        "00100010", -- 0x1F57
        "10101110", -- 0x1F58
        "10000011", -- 0x1F59
        "10101111", -- 0x1F5A
        "10000010", -- 0x1F5B
        "10100011", -- 0x1F5C
        "11100000", -- 0x1F5D
        "00100100", -- 0x1F5E
        "00000001", -- 0x1F5F
        "11110000", -- 0x1F60
        "11001111", -- 0x1F61
        "11110101", -- 0x1F62
        "10000010", -- 0x1F63
        "10001110", -- 0x1F64
        "10000011", -- 0x1F65
        "11100000", -- 0x1F66
        "00110100", -- 0x1F67
        "00000000", -- 0x1F68
        "11110000", -- 0x1F69
        "11111110", -- 0x1F6A
        "00100010", -- 0x1F6B
        "01110101", -- 0x1F6C
        "11100101", -- 0x1F6D
        "00000000", -- 0x1F6E
        "01110101", -- 0x1F6F
        "10110000", -- 0x1F70
        "00000000", -- 0x1F71
        "01010011", -- 0x1F72
        "11010101", -- 0x1F73
        "11110011", -- 0x1F74
        "01000011", -- 0x1F75
        "11010101", -- 0x1F76
        "00001000", -- 0x1F77
        "01010011", -- 0x1F78
        "11010101", -- 0x1F79
        "11001111", -- 0x1F7A
        "01000011", -- 0x1F7B
        "11010101", -- 0x1F7C
        "00100000", -- 0x1F7D
        "00100010", -- 0x1F7E
        "10101000", -- 0x1F7F
        "11101110", -- 0x1F80
        "10001111", -- 0x1F81
        "11111110", -- 0x1F82
        "10001101", -- 0x1F83
        "11110110", -- 0x1F84
        "01110101", -- 0x1F85
        "11101110", -- 0x1F86
        "00000010", -- 0x1F87
        "11100100", -- 0x1F88
        "11111110", -- 0x1F89
        "11111101", -- 0x1F8A
        "11111100", -- 0x1F8B
        "01111111", -- 0x1F8C
        "00000101", -- 0x1F8D
        "00000010", -- 0x1F8E
        "00010110", -- 0x1F8F
        "00110100", -- 0x1F90
        "10100011", -- 0x1F91
        "11100000", -- 0x1F92
        "00101111", -- 0x1F93
        "11111111", -- 0x1F94
        "11110000", -- 0x1F95
        "11100101", -- 0x1F96
        "10000010", -- 0x1F97
        "01110000", -- 0x1F98
        "00000010", -- 0x1F99
        "00010101", -- 0x1F9A
        "10000011", -- 0x1F9B
        "00010101", -- 0x1F9C
        "10000010", -- 0x1F9D
        "11100000", -- 0x1F9E
        "00111110", -- 0x1F9F
        "11111110", -- 0x1FA0
        "11110000", -- 0x1FA1
        "00100010", -- 0x1FA2
        "00010010", -- 0x1FA3
        "00100010", -- 0x1FA4
        "10101100", -- 0x1FA5
        "10010000", -- 0x1FA6
        "00000001", -- 0x1FA7
        "01010001", -- 0x1FA8
        "11100000", -- 0x1FA9
        "00010010", -- 0x1FAA
        "00100100", -- 0x1FAB
        "01000010", -- 0x1FAC
        "00010010", -- 0x1FAD
        "00100100", -- 0x1FAE
        "00010010", -- 0x1FAF
        "01111111", -- 0x1FB0
        "00001100", -- 0x1FB1
        "00000010", -- 0x1FB2
        "00010001", -- 0x1FB3
        "11110101", -- 0x1FB4
        "10010000", -- 0x1FB5
        "00000000", -- 0x1FB6
        "00000001", -- 0x1FB7
        "11100100", -- 0x1FB8
        "11110000", -- 0x1FB9
        "10001111", -- 0x1FBA
        "11111111", -- 0x1FBB
        "10000000", -- 0x1FBC
        "00000001", -- 0x1FBD
        "00000000", -- 0x1FBE
        "10010000", -- 0x1FBF
        "00000000", -- 0x1FC0
        "00000001", -- 0x1FC1
        "11100000", -- 0x1FC2
        "01100000", -- 0x1FC3
        "11111001", -- 0x1FC4
        "00100010", -- 0x1FC5
        "00010010", -- 0x1FC6
        "00100100", -- 0x1FC7
        "10000111", -- 0x1FC8
        "00101000", -- 0x1FC9
        "11111001", -- 0x1FCA
        "11100100", -- 0x1FCB
        "00110011", -- 0x1FCC
        "11111000", -- 0x1FCD
        "10100011", -- 0x1FCE
        "11100000", -- 0x1FCF
        "11111010", -- 0x1FD0
        "00101001", -- 0x1FD1
        "11111001", -- 0x1FD2
        "11100100", -- 0x1FD3
        "00111000", -- 0x1FD4
        "11111000", -- 0x1FD5
        "00100010", -- 0x1FD6
        "11111111", -- 0x1FD7
        "01111101", -- 0x1FD8
        "00000010", -- 0x1FD9
        "01111110", -- 0x1FDA
        "00000000", -- 0x1FDB
        "00010010", -- 0x1FDC
        "00100000", -- 0x1FDD
        "00001001", -- 0x1FDE
        "11101111", -- 0x1FDF
        "00100100", -- 0x1FE0
        "00001001", -- 0x1FE1
        "11111111", -- 0x1FE2
        "11101110", -- 0x1FE3
        "00110100", -- 0x1FE4
        "00000010", -- 0x1FE5
        "11111110", -- 0x1FE6
        "00100010", -- 0x1FE7
        "00000101", -- 0x1FE8
        "00000001", -- 0x1FE9
        "00000000", -- 0x1FEA
        "00000000", -- 0x1FEB
        "00000000", -- 0x1FEC
        "00110111", -- 0x1FED
        "00000001", -- 0x1FEE
        "00011000", -- 0x1FEF
        "00000101", -- 0x1FF0
        "00000010", -- 0x1FF1
        "00000001", -- 0x1FF2
        "00011000", -- 0x1FF3
        "00000000", -- 0x1FF4
        "00000000", -- 0x1FF5
        "00010110", -- 0x1FF6
        "10111000", -- 0x1FF7
        "00000000", -- 0x1FF8
        "11100101", -- 0x1FF9
        "00001100", -- 0x1FFA
        "00100100", -- 0x1FFB
        "00000011", -- 0x1FFC
        "11111011", -- 0x1FFD
        "11100100", -- 0x1FFE
        "00110101", -- 0x1FFF
        "00001011", -- 0x2000
        "11111010", -- 0x2001
        "10001011", -- 0x2002
        "10000010", -- 0x2003
        "10001010", -- 0x2004
        "10000011", -- 0x2005
        "11100000", -- 0x2006
        "11111001", -- 0x2007
        "00100010", -- 0x2008
        "11101101", -- 0x2009
        "01010100", -- 0x200A
        "00001111", -- 0x200B
        "01100000", -- 0x200C
        "00001010", -- 0x200D
        "11111101", -- 0x200E
        "11101111", -- 0x200F
        "00100101", -- 0x2010
        "11100000", -- 0x2011
        "11001110", -- 0x2012
        "00110011", -- 0x2013
        "11001110", -- 0x2014
        "11011101", -- 0x2015
        "11111001", -- 0x2016
        "11111111", -- 0x2017
        "00100010", -- 0x2018
        "11101101", -- 0x2019
        "01010100", -- 0x201A
        "00001111", -- 0x201B
        "01100000", -- 0x201C
        "00001010", -- 0x201D
        "11111101", -- 0x201E
        "11101110", -- 0x201F
        "11000011", -- 0x2020
        "00010011", -- 0x2021
        "11001111", -- 0x2022
        "00010011", -- 0x2023
        "11001111", -- 0x2024
        "11011101", -- 0x2025
        "11111001", -- 0x2026
        "11111110", -- 0x2027
        "00100010", -- 0x2028
        "10010000", -- 0x2029
        "00000000", -- 0x202A
        "00000010", -- 0x202B
        "11100000", -- 0x202C
        "10010000", -- 0x202D
        "00000001", -- 0x202E
        "01100001", -- 0x202F
        "00010010", -- 0x2030
        "00100010", -- 0x2031
        "11101011", -- 0x2032
        "11100000", -- 0x2033
        "10010000", -- 0x2034
        "00011000", -- 0x2035
        "00100000", -- 0x2036
        "11110000", -- 0x2037
        "00100010", -- 0x2038
        "01010100", -- 0x2039
        "00001111", -- 0x203A
        "00010010", -- 0x203B
        "00100011", -- 0x203C
        "01001110", -- 0x203D
        "10010000", -- 0x203E
        "00000001", -- 0x203F
        "01010010", -- 0x2040
        "11101110", -- 0x2041
        "11110000", -- 0x2042
        "11101111", -- 0x2043
        "10100011", -- 0x2044
        "11110000", -- 0x2045
        "00000010", -- 0x2046
        "00100100", -- 0x2047
        "01001000", -- 0x2048
        "10010000", -- 0x2049
        "00000110", -- 0x204A
        "10001010", -- 0x204B
        "11100000", -- 0x204C
        "11111101", -- 0x204D
        "01111100", -- 0x204E
        "00000000", -- 0x204F
        "01111110", -- 0x2050
        "00000000", -- 0x2051
        "01111111", -- 0x2052
        "00001010", -- 0x2053
        "00010010", -- 0x2054
        "00011110", -- 0x2055
        "10110110", -- 0x2056
        "11101111", -- 0x2057
        "00100010", -- 0x2058
        "11100100", -- 0x2059
        "11111110", -- 0x205A
        "11111101", -- 0x205B
        "11111100", -- 0x205C
        "01111111", -- 0x205D
        "00000110", -- 0x205E
        "00010010", -- 0x205F
        "00010110", -- 0x2060
        "00110100", -- 0x2061
        "11100101", -- 0x2062
        "10110101", -- 0x2063
        "11111001", -- 0x2064
        "01111000", -- 0x2065
        "00000000", -- 0x2066
        "00100010", -- 0x2067
        "11100101", -- 0x2068
        "00001100", -- 0x2069
        "00100100", -- 0x206A
        "00000010", -- 0x206B
        "11111001", -- 0x206C
        "11100100", -- 0x206D
        "00110101", -- 0x206E
        "00001011", -- 0x206F
        "00010010", -- 0x2070
        "00100100", -- 0x2071
        "10011001", -- 0x2072
        "11111001", -- 0x2073
        "01111000", -- 0x2074
        "00000000", -- 0x2075
        "00100010", -- 0x2076
        "00010010", -- 0x2077
        "00100010", -- 0x2078
        "10111110", -- 0x2079
        "01110100", -- 0x207A
        "00011100", -- 0x207B
        "11110000", -- 0x207C
        "10100011", -- 0x207D
        "01110100", -- 0x207E
        "00100000", -- 0x207F
        "00010010", -- 0x2080
        "00100011", -- 0x2081
        "00110110", -- 0x2082
        "00000010", -- 0x2083
        "00100100", -- 0x2084
        "00101010", -- 0x2085
        "00010010", -- 0x2086
        "00100011", -- 0x2087
        "11110001", -- 0x2088
        "10010000", -- 0x2089
        "00000001", -- 0x208A
        "01100001", -- 0x208B
        "10001101", -- 0x208C
        "00000111", -- 0x208D
        "10001100", -- 0x208E
        "00000110", -- 0x208F
        "00010010", -- 0x2090
        "00100001", -- 0x2091
        "11101011", -- 0x2092
        "11100000", -- 0x2093
        "00100010", -- 0x2094
        "11111000", -- 0x2095
        "10010000", -- 0x2096
        "00010111", -- 0x2097
        "11011111", -- 0x2098
        "10101101", -- 0x2099
        "00000001", -- 0x209A
        "10101100", -- 0x209B
        "00000000", -- 0x209C
        "01111110", -- 0x209D
        "00000000", -- 0x209E
        "01111111", -- 0x209F
        "00001010", -- 0x20A0
        "00000010", -- 0x20A1
        "00011101", -- 0x20A2
        "10000110", -- 0x20A3
        "10010000", -- 0x20A4
        "00000111", -- 0x20A5
        "11001101", -- 0x20A6
        "11100100", -- 0x20A7
        "11110000", -- 0x20A8
        "10100011", -- 0x20A9
        "10100011", -- 0x20AA
        "11100100", -- 0x20AB
        "11110000", -- 0x20AC
        "10010000", -- 0x20AD
        "00000111", -- 0x20AE
        "11001110", -- 0x20AF
        "11100100", -- 0x20B0
        "11110000", -- 0x20B1
        "00100010", -- 0x20B2
        "00010010", -- 0x20B3
        "00100011", -- 0x20B4
        "00011110", -- 0x20B5
        "01110100", -- 0x20B6
        "00010000", -- 0x20B7
        "00010010", -- 0x20B8
        "00100011", -- 0x20B9
        "10001000", -- 0x20BA
        "10010000", -- 0x20BB
        "00011000", -- 0x20BC
        "00001000", -- 0x20BD
        "01110100", -- 0x20BE
        "00000010", -- 0x20BF
        "00100010", -- 0x20C0
        "11111001", -- 0x20C1
        "11100100", -- 0x20C2
        "00110101", -- 0x20C3
        "00001011", -- 0x20C4
        "00010010", -- 0x20C5
        "00100100", -- 0x20C6
        "10011001", -- 0x20C7
        "00010010", -- 0x20C8
        "00100100", -- 0x20C9
        "01000010", -- 0x20CA
        "10010000", -- 0x20CB
        "00010111", -- 0x20CC
        "11010011", -- 0x20CD
        "00100010", -- 0x20CE
        "10010000", -- 0x20CF
        "00000000", -- 0x20D0
        "00000000", -- 0x20D1
        "11100000", -- 0x20D2
        "11111000", -- 0x20D3
        "10010000", -- 0x20D4
        "00000000", -- 0x20D5
        "00000010", -- 0x20D6
        "11100000", -- 0x20D7
        "11111001", -- 0x20D8
        "11101000", -- 0x20D9
        "11000011", -- 0x20DA
        "10011001", -- 0x20DB
        "00100010", -- 0x20DC
        "11100101", -- 0x20DD
        "11011100", -- 0x20DE
        "00010010", -- 0x20DF
        "00100010", -- 0x20E0
        "01101000", -- 0x20E1
        "11111000", -- 0x20E2
        "11100101", -- 0x20E3
        "11011100", -- 0x20E4
        "00010010", -- 0x20E5
        "00100010", -- 0x20E6
        "01011110", -- 0x20E7
        "11111001", -- 0x20E8
        "00100010", -- 0x20E9
        "00010010", -- 0x20EA
        "00100001", -- 0x20EB
        "11001000", -- 0x20EC
        "11100101", -- 0x20ED
        "11000100", -- 0x20EE
        "00010010", -- 0x20EF
        "00100100", -- 0x20F0
        "01000010", -- 0x20F1
        "01110100", -- 0x20F2
        "00011000", -- 0x20F3
        "00000010", -- 0x20F4
        "00011111", -- 0x20F5
        "00110000", -- 0x20F6
        "00010010", -- 0x20F7
        "00100001", -- 0x20F8
        "11001000", -- 0x20F9
        "11100101", -- 0x20FA
        "10110100", -- 0x20FB
        "00010010", -- 0x20FC
        "00100100", -- 0x20FD
        "01000010", -- 0x20FE
        "01110100", -- 0x20FF
        "00001000", -- 0x2100
        "00000010", -- 0x2101
        "00011111", -- 0x2102
        "00110000", -- 0x2103
        "11100000", -- 0x2104
        "11111000", -- 0x2105
        "01111001", -- 0x2106
        "00000000", -- 0x2107
        "11101001", -- 0x2108
        "00100100", -- 0x2109
        "11010000", -- 0x210A
        "11111111", -- 0x210B
        "11101000", -- 0x210C
        "00110100", -- 0x210D
        "00000111", -- 0x210E
        "11111110", -- 0x210F
        "00100010", -- 0x2110
        "01010100", -- 0x2111
        "00001111", -- 0x2112
        "00010010", -- 0x2113
        "00100011", -- 0x2114
        "01001110", -- 0x2115
        "10010000", -- 0x2116
        "00000001", -- 0x2117
        "01010110", -- 0x2118
        "11101110", -- 0x2119
        "11110000", -- 0x211A
        "11101111", -- 0x211B
        "10100011", -- 0x211C
        "00100010", -- 0x211D
        "10010000", -- 0x211E
        "00011000", -- 0x211F
        "00101101", -- 0x2120
        "00010010", -- 0x2121
        "00100001", -- 0x2122
        "11001000", -- 0x2123
        "11100100", -- 0x2124
        "11111101", -- 0x2125
        "11111100", -- 0x2126
        "10010000", -- 0x2127
        "00011000", -- 0x2128
        "00101101", -- 0x2129
        "00100010", -- 0x212A
        "10010000", -- 0x212B
        "00000001", -- 0x212C
        "01010101", -- 0x212D
        "11100000", -- 0x212E
        "11111101", -- 0x212F
        "00011101", -- 0x2130
        "01111110", -- 0x2131
        "00000000", -- 0x2132
        "01111111", -- 0x2133
        "11001000", -- 0x2134
        "00000010", -- 0x2135
        "00100000", -- 0x2136
        "00001001", -- 0x2137
        "00010010", -- 0x2138
        "00011101", -- 0x2139
        "00110011", -- 0x213A
        "00010010", -- 0x213B
        "00011110", -- 0x213C
        "01110100", -- 0x213D
        "00010010", -- 0x213E
        "00011110", -- 0x213F
        "01011101", -- 0x2140
        "00000010", -- 0x2141
        "00100000", -- 0x2142
        "10100100", -- 0x2143
        "10010000", -- 0x2144
        "00000001", -- 0x2145
        "01010100", -- 0x2146
        "00010010", -- 0x2147
        "00100100", -- 0x2148
        "01110011", -- 0x2149
        "10010000", -- 0x214A
        "00000001", -- 0x214B
        "01010010", -- 0x214C
        "00000010", -- 0x214D
        "00100010", -- 0x214E
        "00001100", -- 0x214F
        "00010010", -- 0x2150
        "00100001", -- 0x2151
        "10111100", -- 0x2152
        "01110100", -- 0x2153
        "00001000", -- 0x2154
        "00010010", -- 0x2155
        "00011111", -- 0x2156
        "00011100", -- 0x2157
        "11101111", -- 0x2158
        "11110101", -- 0x2159
        "11101111", -- 0x215A
        "00100010", -- 0x215B
        "10100100", -- 0x215C
        "00100101", -- 0x215D
        "10000010", -- 0x215E
        "11110101", -- 0x215F
        "10000010", -- 0x2160
        "11100101", -- 0x2161
        "10000011", -- 0x2162
        "00110101", -- 0x2163
        "11110000", -- 0x2164
        "11110101", -- 0x2165
        "10000011", -- 0x2166
        "00100010", -- 0x2167
        "11110000", -- 0x2168
        "11100101", -- 0x2169
        "00001100", -- 0x216A
        "00100100", -- 0x216B
        "00000011", -- 0x216C
        "11111001", -- 0x216D
        "11100100", -- 0x216E
        "00110101", -- 0x216F
        "00001011", -- 0x2170
        "00000010", -- 0x2171
        "00100100", -- 0x2172
        "10011001", -- 0x2173
        "11101100", -- 0x2174
        "11110000", -- 0x2175
        "11101101", -- 0x2176
        "10100011", -- 0x2177
        "11110000", -- 0x2178
        "11101110", -- 0x2179
        "10100011", -- 0x217A
        "11110000", -- 0x217B
        "11101111", -- 0x217C
        "10100011", -- 0x217D
        "11110000", -- 0x217E
        "00100010", -- 0x217F
        "11100000", -- 0x2180
        "11111010", -- 0x2181
        "00101001", -- 0x2182
        "11111111", -- 0x2183
        "11100100", -- 0x2184
        "00111000", -- 0x2185
        "11111110", -- 0x2186
        "01111101", -- 0x2187
        "00000010", -- 0x2188
        "00000010", -- 0x2189
        "00100000", -- 0x218A
        "00011001", -- 0x218B
        "10010000", -- 0x218C
        "00000011", -- 0x218D
        "10000110", -- 0x218E
        "11100000", -- 0x218F
        "11111111", -- 0x2190
        "01111101", -- 0x2191
        "00000010", -- 0x2192
        "01111110", -- 0x2193
        "00000000", -- 0x2194
        "00000010", -- 0x2195
        "00100000", -- 0x2196
        "00001001", -- 0x2197
        "10010000", -- 0x2198
        "00000001", -- 0x2199
        "10110101", -- 0x219A
        "11100000", -- 0x219B
        "11111111", -- 0x219C
        "01111101", -- 0x219D
        "00000011", -- 0x219E
        "01111110", -- 0x219F
        "00000000", -- 0x21A0
        "00000010", -- 0x21A1
        "00100000", -- 0x21A2
        "00001001", -- 0x21A3
        "11000000", -- 0x21A4
        "00000100", -- 0x21A5
        "11000000", -- 0x21A6
        "00000101", -- 0x21A7
        "11000000", -- 0x21A8
        "00000110", -- 0x21A9
        "11000000", -- 0x21AA
        "00000111", -- 0x21AB
        "00010010", -- 0x21AC
        "00011100", -- 0x21AD
        "01000000", -- 0x21AE
        "00100010", -- 0x21AF
        "00010010", -- 0x21B0
        "00100001", -- 0x21B1
        "10011000", -- 0x21B2
        "11100101", -- 0x21B3
        "00010111", -- 0x21B4
        "00101111", -- 0x21B5
        "11111001", -- 0x21B6
        "11100101", -- 0x21B7
        "00010110", -- 0x21B8
        "00111110", -- 0x21B9
        "11111000", -- 0x21BA
        "00100010", -- 0x21BB
        "11100000", -- 0x21BC
        "11111100", -- 0x21BD
        "10100011", -- 0x21BE
        "11100000", -- 0x21BF
        "11111101", -- 0x21C0
        "10100011", -- 0x21C1
        "11100000", -- 0x21C2
        "11111110", -- 0x21C3
        "10100011", -- 0x21C4
        "11100000", -- 0x21C5
        "11111111", -- 0x21C6
        "00100010", -- 0x21C7
        "11101100", -- 0x21C8
        "11110000", -- 0x21C9
        "10100011", -- 0x21CA
        "11101101", -- 0x21CB
        "11110000", -- 0x21CC
        "10100011", -- 0x21CD
        "11101110", -- 0x21CE
        "11110000", -- 0x21CF
        "10100011", -- 0x21D0
        "11101111", -- 0x21D1
        "11110000", -- 0x21D2
        "00100010", -- 0x21D3
        "11110000", -- 0x21D4
        "00010010", -- 0x21D5
        "00100011", -- 0x21D6
        "01110011", -- 0x21D7
        "01110100", -- 0x21D8
        "10100001", -- 0x21D9
        "11110000", -- 0x21DA
        "10100011", -- 0x21DB
        "11100100", -- 0x21DC
        "11110000", -- 0x21DD
        "10100011", -- 0x21DE
        "00100010", -- 0x21DF
        "10010000", -- 0x21E0
        "00000010", -- 0x21E1
        "00001000", -- 0x21E2
        "11100100", -- 0x21E3
        "11110000", -- 0x21E4
        "10010000", -- 0x21E5
        "00000001", -- 0x21E6
        "00011010", -- 0x21E7
        "11100100", -- 0x21E8
        "11110000", -- 0x21E9
        "00100010", -- 0x21EA
        "11101111", -- 0x21EB
        "00100101", -- 0x21EC
        "10000010", -- 0x21ED
        "11110101", -- 0x21EE
        "10000010", -- 0x21EF
        "11101110", -- 0x21F0
        "00110101", -- 0x21F1
        "10000011", -- 0x21F2
        "11110101", -- 0x21F3
        "10000011", -- 0x21F4
        "00100010", -- 0x21F5
        "11100101", -- 0x21F6
        "00001100", -- 0x21F7
        "00100100", -- 0x21F8
        "00000011", -- 0x21F9
        "11111001", -- 0x21FA
        "11100100", -- 0x21FB
        "00110101", -- 0x21FC
        "00001011", -- 0x21FD
        "00000010", -- 0x21FE
        "00100100", -- 0x21FF
        "10011001", -- 0x2200
        "00001111", -- 0x2201
        "10111111", -- 0x2202
        "00000000", -- 0x2203
        "00000001", -- 0x2204
        "00001110", -- 0x2205
        "10001111", -- 0x2206
        "10000010", -- 0x2207
        "10001110", -- 0x2208
        "10000011", -- 0x2209
        "11100000", -- 0x220A
        "00100010", -- 0x220B
        "11100000", -- 0x220C
        "11111010", -- 0x220D
        "10100011", -- 0x220E
        "11100000", -- 0x220F
        "11111011", -- 0x2210
        "11101001", -- 0x2211
        "11000011", -- 0x2212
        "10011011", -- 0x2213
        "11101000", -- 0x2214
        "10011010", -- 0x2215
        "00100010", -- 0x2216
        "01111110", -- 0x2217
        "00000001", -- 0x2218
        "01111111", -- 0x2219
        "10000101", -- 0x221A
        "01111100", -- 0x221B
        "00000000", -- 0x221C
        "01111101", -- 0x221D
        "00110000", -- 0x221E
        "00000010", -- 0x221F
        "00011011", -- 0x2220
        "00110101", -- 0x2221
        "10010000", -- 0x2222
        "00000001", -- 0x2223
        "01011000", -- 0x2224
        "00010010", -- 0x2225
        "00100011", -- 0x2226
        "11010101", -- 0x2227
        "10010000", -- 0x2228
        "00000001", -- 0x2229
        "01010100", -- 0x222A
        "00100010", -- 0x222B
        "10010000", -- 0x222C
        "00000001", -- 0x222D
        "01010100", -- 0x222E
        "00010010", -- 0x222F
        "00100011", -- 0x2230
        "11010101", -- 0x2231
        "10010000", -- 0x2232
        "00000001", -- 0x2233
        "01011000", -- 0x2234
        "00100010", -- 0x2235
        "11110000", -- 0x2236
        "10100011", -- 0x2237
        "11100100", -- 0x2238
        "11110000", -- 0x2239
        "00010010", -- 0x223A
        "00100100", -- 0x223B
        "00110000", -- 0x223C
        "11110000", -- 0x223D
        "10100011", -- 0x223E
        "00100010", -- 0x223F
        "11100101", -- 0x2240
        "10111100", -- 0x2241
        "00010010", -- 0x2242
        "00100100", -- 0x2243
        "01000010", -- 0x2244
        "01110100", -- 0x2245
        "00010000", -- 0x2246
        "00000010", -- 0x2247
        "00011111", -- 0x2248
        "00110000", -- 0x2249
        "11100000", -- 0x224A
        "11111111", -- 0x224B
        "01111110", -- 0x224C
        "00000000", -- 0x224D
        "00001111", -- 0x224E
        "10111111", -- 0x224F
        "00000000", -- 0x2250
        "00000001", -- 0x2251
        "00001110", -- 0x2252
        "00100010", -- 0x2253
        "00010010", -- 0x2254
        "00100011", -- 0x2255
        "11000111", -- 0x2256
        "01010011", -- 0x2257
        "11101101", -- 0x2258
        "11001111", -- 0x2259
        "01000011", -- 0x225A
        "11101101", -- 0x225B
        "00100000", -- 0x225C
        "00100010", -- 0x225D
        "01010100", -- 0x225E
        "11000000", -- 0x225F
        "01100100", -- 0x2260
        "01000000", -- 0x2261
        "00100100", -- 0x2262
        "11111111", -- 0x2263
        "10110011", -- 0x2264
        "11100100", -- 0x2265
        "00110011", -- 0x2266
        "00100010", -- 0x2267
        "01010100", -- 0x2268
        "00110000", -- 0x2269
        "01100100", -- 0x226A
        "00010000", -- 0x226B
        "00100100", -- 0x226C
        "11111111", -- 0x226D
        "10110011", -- 0x226E
        "11100100", -- 0x226F
        "00110011", -- 0x2270
        "00100010", -- 0x2271
        "00010010", -- 0x2272
        "00100011", -- 0x2273
        "01010110", -- 0x2274
        "01111111", -- 0x2275
        "01001100", -- 0x2276
        "00010010", -- 0x2277
        "00010001", -- 0x2278
        "11110101", -- 0x2279
        "11100100", -- 0x227A
        "00100010", -- 0x227B
        "00010010", -- 0x227C
        "00100000", -- 0x227D
        "10110011", -- 0x227E
        "11110000", -- 0x227F
        "10100011", -- 0x2280
        "11100100", -- 0x2281
        "11110000", -- 0x2282
        "00000010", -- 0x2283
        "00100011", -- 0x2284
        "01111010", -- 0x2285
        "11100100", -- 0x2286
        "11111110", -- 0x2287
        "11111101", -- 0x2288
        "11111100", -- 0x2289
        "10010000", -- 0x228A
        "00011000", -- 0x228B
        "00101101", -- 0x228C
        "01111111", -- 0x228D
        "00001010", -- 0x228E
        "00100010", -- 0x228F
        "01110100", -- 0x2290
        "11100001", -- 0x2291
        "11110000", -- 0x2292
        "10100011", -- 0x2293
        "10100011", -- 0x2294
        "11100100", -- 0x2295
        "11110000", -- 0x2296
        "10100011", -- 0x2297
        "11110000", -- 0x2298
        "00100010", -- 0x2299
        "00010010", -- 0x229A
        "00011011", -- 0x229B
        "00001101", -- 0x229C
        "00010010", -- 0x229D
        "00100011", -- 0x229E
        "11100011", -- 0x229F
        "00000010", -- 0x22A0
        "00011111", -- 0x22A1
        "01101100", -- 0x22A2
        "00010010", -- 0x22A3
        "00010111", -- 0x22A4
        "11010001", -- 0x22A5
        "10010000", -- 0x22A6
        "00000100", -- 0x22A7
        "10000111", -- 0x22A8
        "11100100", -- 0x22A9
        "11110000", -- 0x22AA
        "00100010", -- 0x22AB
        "00010010", -- 0x22AC
        "00010101", -- 0x22AD
        "10010000", -- 0x22AE
        "10010000", -- 0x22AF
        "00000011", -- 0x22B0
        "10000111", -- 0x22B1
        "11100100", -- 0x22B2
        "11110000", -- 0x22B3
        "00100010", -- 0x22B4
        "01111111", -- 0x22B5
        "00001000", -- 0x22B6
        "00010010", -- 0x22B7
        "00011110", -- 0x22B8
        "10001011", -- 0x22B9
        "11100101", -- 0x22BA
        "10101101", -- 0x22BB
        "11111111", -- 0x22BC
        "00100010", -- 0x22BD
        "11110000", -- 0x22BE
        "00010010", -- 0x22BF
        "00100011", -- 0x22C0
        "01110011", -- 0x22C1
        "01110100", -- 0x22C2
        "00001001", -- 0x22C3
        "11110000", -- 0x22C4
        "10100011", -- 0x22C5
        "00100010", -- 0x22C6
        "11110000", -- 0x22C7
        "00010010", -- 0x22C8
        "00100011", -- 0x22C9
        "01110011", -- 0x22CA
        "01110100", -- 0x22CB
        "00000001", -- 0x22CC
        "11110000", -- 0x22CD
        "10100011", -- 0x22CE
        "00100010", -- 0x22CF
        "11110000", -- 0x22D0
        "00010010", -- 0x22D1
        "00100011", -- 0x22D2
        "01110011", -- 0x22D3
        "01110100", -- 0x22D4
        "10100000", -- 0x22D5
        "11110000", -- 0x22D6
        "10100011", -- 0x22D7
        "00100010", -- 0x22D8
        "11111011", -- 0x22D9
        "11100100", -- 0x22DA
        "00111000", -- 0x22DB
        "11111010", -- 0x22DC
        "10001011", -- 0x22DD
        "10000010", -- 0x22DE
        "10001010", -- 0x22DF
        "10000011", -- 0x22E0
        "00100010", -- 0x22E1
        "01111100", -- 0x22E2
        "00000001", -- 0x22E3
        "01111101", -- 0x22E4
        "00000000", -- 0x22E5
        "01111110", -- 0x22E6
        "00000101", -- 0x22E7
        "01111111", -- 0x22E8
        "10001001", -- 0x22E9
        "00100010", -- 0x22EA
        "00100101", -- 0x22EB
        "10000010", -- 0x22EC
        "11110101", -- 0x22ED
        "10000010", -- 0x22EE
        "01010000", -- 0x22EF
        "00000010", -- 0x22F0
        "00000101", -- 0x22F1
        "10000011", -- 0x22F2
        "00100010", -- 0x22F3
        "10010000", -- 0x22F4
        "00000110", -- 0x22F5
        "10001010", -- 0x22F6
        "11100000", -- 0x22F7
        "00000100", -- 0x22F8
        "01010100", -- 0x22F9
        "00011111", -- 0x22FA
        "11110000", -- 0x22FB
        "00100010", -- 0x22FC
        "10010000", -- 0x22FD
        "00000001", -- 0x22FE
        "10010011", -- 0x22FF
        "11100000", -- 0x2300
        "11111010", -- 0x2301
        "10100011", -- 0x2302
        "11100000", -- 0x2303
        "11111011", -- 0x2304
        "00100010", -- 0x2305
        "10000101", -- 0x2306
        "00001100", -- 0x2307
        "10000010", -- 0x2308
        "10000101", -- 0x2309
        "00001011", -- 0x230A
        "10000011", -- 0x230B
        "11100000", -- 0x230C
        "00100010", -- 0x230D
        "11110000", -- 0x230E
        "00010010", -- 0x230F
        "00100011", -- 0x2310
        "01110011", -- 0x2311
        "01110100", -- 0x2312
        "00000110", -- 0x2313
        "11110000", -- 0x2314
        "00100010", -- 0x2315
        "00010010", -- 0x2316
        "00100011", -- 0x2317
        "10011101", -- 0x2318
        "01110100", -- 0x2319
        "00000001", -- 0x231A
        "00000010", -- 0x231B
        "00100100", -- 0x231C
        "01011010", -- 0x231D
        "10010000", -- 0x231E
        "00011000", -- 0x231F
        "00000111", -- 0x2320
        "01110100", -- 0x2321
        "00010101", -- 0x2322
        "11110000", -- 0x2323
        "10100011", -- 0x2324
        "00100010", -- 0x2325
        "00010010", -- 0x2326
        "00100001", -- 0x2327
        "11001000", -- 0x2328
        "11100101", -- 0x2329
        "10101100", -- 0x232A
        "00000010", -- 0x232B
        "00100100", -- 0x232C
        "01000010", -- 0x232D
        "10010000", -- 0x232E
        "00000001", -- 0x232F
        "00101001", -- 0x2330
        "11100100", -- 0x2331
        "11111110", -- 0x2332
        "11111101", -- 0x2333
        "11111100", -- 0x2334
        "00100010", -- 0x2335
        "00010010", -- 0x2336
        "00100011", -- 0x2337
        "10001111", -- 0x2338
        "11110000", -- 0x2339
        "10100011", -- 0x233A
        "11100100", -- 0x233B
        "11110000", -- 0x233C
        "00100010", -- 0x233D
        "11111001", -- 0x233E
        "11100100", -- 0x233F
        "00110101", -- 0x2340
        "00001111", -- 0x2341
        "11111000", -- 0x2342
        "00000010", -- 0x2343
        "00100100", -- 0x2344
        "10000010", -- 0x2345
        "11100000", -- 0x2346
        "11111110", -- 0x2347
        "10100011", -- 0x2348
        "11100000", -- 0x2349
        "11111111", -- 0x234A
        "00000010", -- 0x234B
        "00100100", -- 0x234C
        "10010101", -- 0x234D
        "11111101", -- 0x234E
        "01111110", -- 0x234F
        "00000000", -- 0x2350
        "01111111", -- 0x2351
        "00000001", -- 0x2352
        "00000010", -- 0x2353
        "00100000", -- 0x2354
        "00001001", -- 0x2355
        "11100100", -- 0x2356
        "11111111", -- 0x2357
        "11111110", -- 0x2358
        "11111101", -- 0x2359
        "11111100", -- 0x235A
        "00000010", -- 0x235B
        "00100100", -- 0x235C
        "00010010", -- 0x235D
        "01111110", -- 0x235E
        "00000011", -- 0x235F
        "01111111", -- 0x2360
        "00101010", -- 0x2361
        "00000010", -- 0x2362
        "00010100", -- 0x2363
        "00010100", -- 0x2364
        "01111110", -- 0x2365
        "00011000", -- 0x2366
        "01111111", -- 0x2367
        "00000111", -- 0x2368
        "00000010", -- 0x2369
        "00010010", -- 0x236A
        "01100111", -- 0x236B
        "01111110", -- 0x236C
        "00000100", -- 0x236D
        "01111111", -- 0x236E
        "11001101", -- 0x236F
        "00000010", -- 0x2370
        "00010100", -- 0x2371
        "00010100", -- 0x2372
        "00010010", -- 0x2373
        "00100011", -- 0x2374
        "01100101", -- 0x2375
        "10010000", -- 0x2376
        "00011000", -- 0x2377
        "00001000", -- 0x2378
        "00100010", -- 0x2379
        "00010010", -- 0x237A
        "00100100", -- 0x237B
        "10010001", -- 0x237C
        "10010000", -- 0x237D
        "00011000", -- 0x237E
        "00001000", -- 0x237F
        "00100010", -- 0x2380
        "11110000", -- 0x2381
        "00010010", -- 0x2382
        "00100011", -- 0x2383
        "01100101", -- 0x2384
        "00000010", -- 0x2385
        "00100011", -- 0x2386
        "00011110", -- 0x2387
        "11110000", -- 0x2388
        "00010010", -- 0x2389
        "00100011", -- 0x238A
        "11001110", -- 0x238B
        "00000010", -- 0x238C
        "00100100", -- 0x238D
        "10001100", -- 0x238E
        "11110000", -- 0x238F
        "00010010", -- 0x2390
        "00100011", -- 0x2391
        "01110011", -- 0x2392
        "01110100", -- 0x2393
        "00001101", -- 0x2394
        "00100010", -- 0x2395
        "11110000", -- 0x2396
        "00010010", -- 0x2397
        "00100100", -- 0x2398
        "00110110", -- 0x2399
        "11110000", -- 0x239A
        "10100011", -- 0x239B
        "00100010", -- 0x239C
        "00010010", -- 0x239D
        "00100010", -- 0x239E
        "11000111", -- 0x239F
        "00010100", -- 0x23A0
        "11110000", -- 0x23A1
        "10100011", -- 0x23A2
        "00100010", -- 0x23A3
        "00010010", -- 0x23A4
        "00011100", -- 0x23A5
        "10001000", -- 0x23A6
        "01001101", -- 0x23A7
        "01001110", -- 0x23A8
        "01001111", -- 0x23A9
        "00100010", -- 0x23AA
        "00010010", -- 0x23AB
        "00011010", -- 0x23AC
        "11100100", -- 0x23AD
        "01001101", -- 0x23AE
        "01001110", -- 0x23AF
        "01001111", -- 0x23B0
        "00100010", -- 0x23B1
        "10010000", -- 0x23B2
        "00000000", -- 0x23B3
        "00000010", -- 0x23B4
        "11100000", -- 0x23B5
        "01111000", -- 0x23B6
        "00000000", -- 0x23B7
        "00100010", -- 0x23B8
        "00010010", -- 0x23B9
        "00010001", -- 0x23BA
        "00000010", -- 0x23BB
        "11100100", -- 0x23BC
        "11111101", -- 0x23BD
        "11111100", -- 0x23BE
        "00100010", -- 0x23BF
        "11101110", -- 0x23C0
        "00110011", -- 0x23C1
        "10010101", -- 0x23C2
        "11100000", -- 0x23C3
        "11111101", -- 0x23C4
        "11111100", -- 0x23C5
        "00100010", -- 0x23C6
        "01010011", -- 0x23C7
        "11101101", -- 0x23C8
        "00111111", -- 0x23C9
        "01000011", -- 0x23CA
        "11101101", -- 0x23CB
        "10000000", -- 0x23CC
        "00100010", -- 0x23CD
        "10100011", -- 0x23CE
        "11100100", -- 0x23CF
        "11110000", -- 0x23D0
        "10010000", -- 0x23D1
        "00011000", -- 0x23D2
        "00001010", -- 0x23D3
        "00100010", -- 0x23D4
        "11100100", -- 0x23D5
        "11110000", -- 0x23D6
        "01110100", -- 0x23D7
        "00000001", -- 0x23D8
        "10100011", -- 0x23D9
        "11110000", -- 0x23DA
        "00100010", -- 0x23DB
        "00100100", -- 0x23DC
        "00000010", -- 0x23DD
        "00010010", -- 0x23DE
        "00100010", -- 0x23DF
        "11011001", -- 0x23E0
        "11100000", -- 0x23E1
        "00100010", -- 0x23E2
        "01110101", -- 0x23E3
        "11111101", -- 0x23E4
        "00010011", -- 0x23E5
        "01110101", -- 0x23E6
        "11110101", -- 0x23E7
        "00010010", -- 0x23E8
        "00100010", -- 0x23E9
        "11111001", -- 0x23EA
        "11100100", -- 0x23EB
        "00111000", -- 0x23EC
        "11111000", -- 0x23ED
        "00000010", -- 0x23EE
        "00100100", -- 0x23EF
        "10000010", -- 0x23F0
        "01111100", -- 0x23F1
        "00000000", -- 0x23F2
        "01111101", -- 0x23F3
        "00100100", -- 0x23F4
        "00000010", -- 0x23F5
        "00010101", -- 0x23F6
        "00110111", -- 0x23F7
        "01111100", -- 0x23F8
        "00000000", -- 0x23F9
        "01111101", -- 0x23FA
        "11001000", -- 0x23FB
        "00000010", -- 0x23FC
        "00100011", -- 0x23FD
        "01101100", -- 0x23FE
        "10001111", -- 0x23FF
        "00000101", -- 0x2400
        "10001110", -- 0x2401
        "00000100", -- 0x2402
        "00000010", -- 0x2403
        "00100011", -- 0x2404
        "01101100", -- 0x2405
        "00010010", -- 0x2406
        "00100011", -- 0x2407
        "00110110", -- 0x2408
        "00000010", -- 0x2409
        "00100011", -- 0x240A
        "01111010", -- 0x240B
        "10010000", -- 0x240C
        "00000001", -- 0x240D
        "01011000", -- 0x240E
        "00000010", -- 0x240F
        "00100100", -- 0x2410
        "10000111", -- 0x2411
        "10010000", -- 0x2412
        "00010111", -- 0x2413
        "11101001", -- 0x2414
        "00000010", -- 0x2415
        "00100001", -- 0x2416
        "11001000", -- 0x2417
        "00010010", -- 0x2418
        "00100100", -- 0x2419
        "01001000", -- 0x241A
        "00000010", -- 0x241B
        "00100100", -- 0x241C
        "01000010", -- 0x241D
        "00010010", -- 0x241E
        "00100011", -- 0x241F
        "10110010", -- 0x2420
        "00100100", -- 0x2421
        "00000011", -- 0x2422
        "00100010", -- 0x2423
        "00010010", -- 0x2424
        "00100100", -- 0x2425
        "01101001", -- 0x2426
        "01100100", -- 0x2427
        "00000001", -- 0x2428
        "00100010", -- 0x2429
        "00010010", -- 0x242A
        "00100100", -- 0x242B
        "10010001", -- 0x242C
        "01111000", -- 0x242D
        "00000000", -- 0x242E
        "00100010", -- 0x242F
        "00010010", -- 0x2430
        "00100011", -- 0x2431
        "01111010", -- 0x2432
        "01110100", -- 0x2433
        "10100001", -- 0x2434
        "00100010", -- 0x2435
        "00010010", -- 0x2436
        "00100011", -- 0x2437
        "01110011", -- 0x2438
        "01110100", -- 0x2439
        "10100010", -- 0x243A
        "00100010", -- 0x243B
        "10010000", -- 0x243C
        "00000001", -- 0x243D
        "10110101", -- 0x243E
        "11100100", -- 0x243F
        "11110000", -- 0x2440
        "00100010", -- 0x2441
        "11111111", -- 0x2442
        "11100100", -- 0x2443
        "11111110", -- 0x2444
        "11111101", -- 0x2445
        "11111100", -- 0x2446
        "00100010", -- 0x2447
        "10001001", -- 0x2448
        "10000010", -- 0x2449
        "10001000", -- 0x244A
        "10000011", -- 0x244B
        "11100000", -- 0x244C
        "00100010", -- 0x244D
        "11100100", -- 0x244E
        "11111101", -- 0x244F
        "11111100", -- 0x2450
        "00000010", -- 0x2451
        "00100011", -- 0x2452
        "01101100", -- 0x2453
        "11101000", -- 0x2454
        "11110000", -- 0x2455
        "11101001", -- 0x2456
        "10100011", -- 0x2457
        "11110000", -- 0x2458
        "00100010", -- 0x2459
        "00010010", -- 0x245A
        "00100011", -- 0x245B
        "00001110", -- 0x245C
        "10100011", -- 0x245D
        "00100010", -- 0x245E
        "00010010", -- 0x245F
        "00100010", -- 0x2460
        "11000111", -- 0x2461
        "10100011", -- 0x2462
        "00100010", -- 0x2463
        "00010010", -- 0x2464
        "00100011", -- 0x2465
        "10010110", -- 0x2466
        "10100011", -- 0x2467
        "00100010", -- 0x2468
        "10010000", -- 0x2469
        "00000001", -- 0x246A
        "00011100", -- 0x246B
        "11100000", -- 0x246C
        "00100010", -- 0x246D
        "10010000", -- 0x246E
        "00000110", -- 0x246F
        "10001001", -- 0x2470
        "11100000", -- 0x2471
        "00100010", -- 0x2472
        "00010010", -- 0x2473
        "00100100", -- 0x2474
        "10000111", -- 0x2475
        "11111001", -- 0x2476
        "00100010", -- 0x2477
        "01010100", -- 0x2478
        "00000111", -- 0x2479
        "00000010", -- 0x247A
        "00100011", -- 0x247B
        "01001110", -- 0x247C
        "01110100", -- 0x247D
        "00000010", -- 0x247E
        "00000010", -- 0x247F
        "00100011", -- 0x2480
        "10001000", -- 0x2481
        "10001001", -- 0x2482
        "10000010", -- 0x2483
        "10001000", -- 0x2484
        "10000011", -- 0x2485
        "00100010", -- 0x2486
        "11100000", -- 0x2487
        "11111000", -- 0x2488
        "10100011", -- 0x2489
        "11100000", -- 0x248A
        "00100010", -- 0x248B
        "11100100", -- 0x248C
        "11110000", -- 0x248D
        "00000010", -- 0x248E
        "00100011", -- 0x248F
        "01100101", -- 0x2490
        "10100011", -- 0x2491
        "00000010", -- 0x2492
        "00100100", -- 0x2493
        "10001100", -- 0x2494
        "11100100", -- 0x2495
        "11111101", -- 0x2496
        "11111100", -- 0x2497
        "00100010", -- 0x2498
        "11111000", -- 0x2499
        "00000010", -- 0x249A
        "00100100", -- 0x249B
        "01001000", -- 0x249C
        "00000010", -- 0x249D
        "00100001", -- 0x249E
        "11100000", -- 0x249F
        "10000000", -- 0x24A0
        "11111110", -- 0x24A1
        "11100100", -- 0x24A2
        "01110011", -- 0x24A3
        "--------", -- 0x24A4
        "--------", -- 0x24A5
        "--------", -- 0x24A6
        "--------", -- 0x24A7
        "--------", -- 0x24A8
        "--------", -- 0x24A9
        "--------", -- 0x24AA
        "--------", -- 0x24AB
        "--------", -- 0x24AC
        "--------", -- 0x24AD
        "--------", -- 0x24AE
        "--------", -- 0x24AF
        "--------", -- 0x24B0
        "--------", -- 0x24B1
        "--------", -- 0x24B2
        "--------", -- 0x24B3
        "--------", -- 0x24B4
        "--------", -- 0x24B5
        "--------", -- 0x24B6
        "--------", -- 0x24B7
        "--------", -- 0x24B8
        "--------", -- 0x24B9
        "--------", -- 0x24BA
        "--------", -- 0x24BB
        "--------", -- 0x24BC
        "--------", -- 0x24BD
        "--------", -- 0x24BE
        "--------", -- 0x24BF
        "--------", -- 0x24C0
        "--------", -- 0x24C1
        "--------", -- 0x24C2
        "--------", -- 0x24C3
        "--------", -- 0x24C4
        "--------", -- 0x24C5
        "--------", -- 0x24C6
        "--------", -- 0x24C7
        "--------", -- 0x24C8
        "--------", -- 0x24C9
        "--------", -- 0x24CA
        "--------", -- 0x24CB
        "--------", -- 0x24CC
        "--------", -- 0x24CD
        "--------", -- 0x24CE
        "--------", -- 0x24CF
        "--------", -- 0x24D0
        "--------", -- 0x24D1
        "--------", -- 0x24D2
        "--------", -- 0x24D3
        "--------", -- 0x24D4
        "--------", -- 0x24D5
        "--------", -- 0x24D6
        "--------", -- 0x24D7
        "--------", -- 0x24D8
        "--------", -- 0x24D9
        "--------", -- 0x24DA
        "--------", -- 0x24DB
        "--------", -- 0x24DC
        "--------", -- 0x24DD
        "--------", -- 0x24DE
        "--------", -- 0x24DF
        "--------", -- 0x24E0
        "--------", -- 0x24E1
        "--------", -- 0x24E2
        "--------", -- 0x24E3
        "--------", -- 0x24E4
        "--------", -- 0x24E5
        "--------", -- 0x24E6
        "--------", -- 0x24E7
        "--------", -- 0x24E8
        "--------", -- 0x24E9
        "--------", -- 0x24EA
        "--------", -- 0x24EB
        "--------", -- 0x24EC
        "--------", -- 0x24ED
        "--------", -- 0x24EE
        "--------", -- 0x24EF
        "--------", -- 0x24F0
        "--------", -- 0x24F1
        "--------", -- 0x24F2
        "--------", -- 0x24F3
        "--------", -- 0x24F4
        "--------", -- 0x24F5
        "--------", -- 0x24F6
        "--------", -- 0x24F7
        "--------", -- 0x24F8
        "--------", -- 0x24F9
        "--------", -- 0x24FA
        "--------", -- 0x24FB
        "--------", -- 0x24FC
        "--------", -- 0x24FD
        "--------", -- 0x24FE
        "--------", -- 0x24FF
        "--------", -- 0x2500
        "--------", -- 0x2501
        "--------", -- 0x2502
        "--------", -- 0x2503
        "--------", -- 0x2504
        "--------", -- 0x2505
        "--------", -- 0x2506
        "--------", -- 0x2507
        "--------", -- 0x2508
        "--------", -- 0x2509
        "--------", -- 0x250A
        "--------", -- 0x250B
        "--------", -- 0x250C
        "--------", -- 0x250D
        "--------", -- 0x250E
        "--------", -- 0x250F
        "--------", -- 0x2510
        "--------", -- 0x2511
        "--------", -- 0x2512
        "--------", -- 0x2513
        "--------", -- 0x2514
        "--------", -- 0x2515
        "--------", -- 0x2516
        "--------", -- 0x2517
        "--------", -- 0x2518
        "--------", -- 0x2519
        "--------", -- 0x251A
        "--------", -- 0x251B
        "--------", -- 0x251C
        "--------", -- 0x251D
        "--------", -- 0x251E
        "--------", -- 0x251F
        "--------", -- 0x2520
        "--------", -- 0x2521
        "--------", -- 0x2522
        "--------", -- 0x2523
        "--------", -- 0x2524
        "--------", -- 0x2525
        "--------", -- 0x2526
        "--------", -- 0x2527
        "--------", -- 0x2528
        "--------", -- 0x2529
        "--------", -- 0x252A
        "--------", -- 0x252B
        "--------", -- 0x252C
        "--------", -- 0x252D
        "--------", -- 0x252E
        "--------", -- 0x252F
        "--------", -- 0x2530
        "--------", -- 0x2531
        "--------", -- 0x2532
        "--------", -- 0x2533
        "--------", -- 0x2534
        "--------", -- 0x2535
        "--------", -- 0x2536
        "--------", -- 0x2537
        "--------", -- 0x2538
        "--------", -- 0x2539
        "--------", -- 0x253A
        "--------", -- 0x253B
        "--------", -- 0x253C
        "--------", -- 0x253D
        "--------", -- 0x253E
        "--------", -- 0x253F
        "--------", -- 0x2540
        "--------", -- 0x2541
        "--------", -- 0x2542
        "--------", -- 0x2543
        "--------", -- 0x2544
        "--------", -- 0x2545
        "--------", -- 0x2546
        "--------", -- 0x2547
        "--------", -- 0x2548
        "--------", -- 0x2549
        "--------", -- 0x254A
        "--------", -- 0x254B
        "--------", -- 0x254C
        "--------", -- 0x254D
        "--------", -- 0x254E
        "--------", -- 0x254F
        "--------", -- 0x2550
        "--------", -- 0x2551
        "--------", -- 0x2552
        "--------", -- 0x2553
        "--------", -- 0x2554
        "--------", -- 0x2555
        "--------", -- 0x2556
        "--------", -- 0x2557
        "--------", -- 0x2558
        "--------", -- 0x2559
        "--------", -- 0x255A
        "--------", -- 0x255B
        "--------", -- 0x255C
        "--------", -- 0x255D
        "--------", -- 0x255E
        "--------", -- 0x255F
        "--------", -- 0x2560
        "--------", -- 0x2561
        "--------", -- 0x2562
        "--------", -- 0x2563
        "--------", -- 0x2564
        "--------", -- 0x2565
        "--------", -- 0x2566
        "--------", -- 0x2567
        "--------", -- 0x2568
        "--------", -- 0x2569
        "--------", -- 0x256A
        "--------", -- 0x256B
        "--------", -- 0x256C
        "--------", -- 0x256D
        "--------", -- 0x256E
        "--------", -- 0x256F
        "--------", -- 0x2570
        "--------", -- 0x2571
        "--------", -- 0x2572
        "--------", -- 0x2573
        "--------", -- 0x2574
        "--------", -- 0x2575
        "--------", -- 0x2576
        "--------", -- 0x2577
        "--------", -- 0x2578
        "--------", -- 0x2579
        "--------", -- 0x257A
        "--------", -- 0x257B
        "--------", -- 0x257C
        "--------", -- 0x257D
        "--------", -- 0x257E
        "--------", -- 0x257F
        "--------", -- 0x2580
        "--------", -- 0x2581
        "--------", -- 0x2582
        "--------", -- 0x2583
        "--------", -- 0x2584
        "--------", -- 0x2585
        "--------", -- 0x2586
        "--------", -- 0x2587
        "--------", -- 0x2588
        "--------", -- 0x2589
        "--------", -- 0x258A
        "--------", -- 0x258B
        "--------", -- 0x258C
        "--------", -- 0x258D
        "--------", -- 0x258E
        "--------", -- 0x258F
        "--------", -- 0x2590
        "--------", -- 0x2591
        "--------", -- 0x2592
        "--------", -- 0x2593
        "--------", -- 0x2594
        "--------", -- 0x2595
        "--------", -- 0x2596
        "--------", -- 0x2597
        "--------", -- 0x2598
        "--------", -- 0x2599
        "--------", -- 0x259A
        "--------", -- 0x259B
        "--------", -- 0x259C
        "--------", -- 0x259D
        "--------", -- 0x259E
        "--------", -- 0x259F
        "--------", -- 0x25A0
        "--------", -- 0x25A1
        "--------", -- 0x25A2
        "--------", -- 0x25A3
        "--------", -- 0x25A4
        "--------", -- 0x25A5
        "--------", -- 0x25A6
        "--------", -- 0x25A7
        "--------", -- 0x25A8
        "--------", -- 0x25A9
        "--------", -- 0x25AA
        "--------", -- 0x25AB
        "--------", -- 0x25AC
        "--------", -- 0x25AD
        "--------", -- 0x25AE
        "--------", -- 0x25AF
        "--------", -- 0x25B0
        "--------", -- 0x25B1
        "--------", -- 0x25B2
        "--------", -- 0x25B3
        "--------", -- 0x25B4
        "--------", -- 0x25B5
        "--------", -- 0x25B6
        "--------", -- 0x25B7
        "--------", -- 0x25B8
        "--------", -- 0x25B9
        "--------", -- 0x25BA
        "--------", -- 0x25BB
        "--------", -- 0x25BC
        "--------", -- 0x25BD
        "--------", -- 0x25BE
        "--------", -- 0x25BF
        "--------", -- 0x25C0
        "--------", -- 0x25C1
        "--------", -- 0x25C2
        "--------", -- 0x25C3
        "--------", -- 0x25C4
        "--------", -- 0x25C5
        "--------", -- 0x25C6
        "--------", -- 0x25C7
        "--------", -- 0x25C8
        "--------", -- 0x25C9
        "--------", -- 0x25CA
        "--------", -- 0x25CB
        "--------", -- 0x25CC
        "--------", -- 0x25CD
        "--------", -- 0x25CE
        "--------", -- 0x25CF
        "--------", -- 0x25D0
        "--------", -- 0x25D1
        "--------", -- 0x25D2
        "--------", -- 0x25D3
        "--------", -- 0x25D4
        "--------", -- 0x25D5
        "--------", -- 0x25D6
        "--------", -- 0x25D7
        "--------", -- 0x25D8
        "--------", -- 0x25D9
        "--------", -- 0x25DA
        "--------", -- 0x25DB
        "--------", -- 0x25DC
        "--------", -- 0x25DD
        "--------", -- 0x25DE
        "--------", -- 0x25DF
        "--------", -- 0x25E0
        "--------", -- 0x25E1
        "--------", -- 0x25E2
        "--------", -- 0x25E3
        "--------", -- 0x25E4
        "--------", -- 0x25E5
        "--------", -- 0x25E6
        "--------", -- 0x25E7
        "--------", -- 0x25E8
        "--------", -- 0x25E9
        "--------", -- 0x25EA
        "--------", -- 0x25EB
        "--------", -- 0x25EC
        "--------", -- 0x25ED
        "--------", -- 0x25EE
        "--------", -- 0x25EF
        "--------", -- 0x25F0
        "--------", -- 0x25F1
        "--------", -- 0x25F2
        "--------", -- 0x25F3
        "--------", -- 0x25F4
        "--------", -- 0x25F5
        "--------", -- 0x25F6
        "--------", -- 0x25F7
        "--------", -- 0x25F8
        "--------", -- 0x25F9
        "--------", -- 0x25FA
        "--------", -- 0x25FB
        "--------", -- 0x25FC
        "--------", -- 0x25FD
        "--------", -- 0x25FE
        "--------", -- 0x25FF
        "--------", -- 0x2600
        "--------", -- 0x2601
        "--------", -- 0x2602
        "--------", -- 0x2603
        "--------", -- 0x2604
        "--------", -- 0x2605
        "--------", -- 0x2606
        "--------", -- 0x2607
        "--------", -- 0x2608
        "--------", -- 0x2609
        "--------", -- 0x260A
        "--------", -- 0x260B
        "--------", -- 0x260C
        "--------", -- 0x260D
        "--------", -- 0x260E
        "--------", -- 0x260F
        "--------", -- 0x2610
        "--------", -- 0x2611
        "--------", -- 0x2612
        "--------", -- 0x2613
        "--------", -- 0x2614
        "--------", -- 0x2615
        "--------", -- 0x2616
        "--------", -- 0x2617
        "--------", -- 0x2618
        "--------", -- 0x2619
        "--------", -- 0x261A
        "--------", -- 0x261B
        "--------", -- 0x261C
        "--------", -- 0x261D
        "--------", -- 0x261E
        "--------", -- 0x261F
        "--------", -- 0x2620
        "--------", -- 0x2621
        "--------", -- 0x2622
        "--------", -- 0x2623
        "--------", -- 0x2624
        "--------", -- 0x2625
        "--------", -- 0x2626
        "--------", -- 0x2627
        "--------", -- 0x2628
        "--------", -- 0x2629
        "--------", -- 0x262A
        "--------", -- 0x262B
        "--------", -- 0x262C
        "--------", -- 0x262D
        "--------", -- 0x262E
        "--------", -- 0x262F
        "--------", -- 0x2630
        "--------", -- 0x2631
        "--------", -- 0x2632
        "--------", -- 0x2633
        "--------", -- 0x2634
        "--------", -- 0x2635
        "--------", -- 0x2636
        "--------", -- 0x2637
        "--------", -- 0x2638
        "--------", -- 0x2639
        "--------", -- 0x263A
        "--------", -- 0x263B
        "--------", -- 0x263C
        "--------", -- 0x263D
        "--------", -- 0x263E
        "--------", -- 0x263F
        "--------", -- 0x2640
        "--------", -- 0x2641
        "--------", -- 0x2642
        "--------", -- 0x2643
        "--------", -- 0x2644
        "--------", -- 0x2645
        "--------", -- 0x2646
        "--------", -- 0x2647
        "--------", -- 0x2648
        "--------", -- 0x2649
        "--------", -- 0x264A
        "--------", -- 0x264B
        "--------", -- 0x264C
        "--------", -- 0x264D
        "--------", -- 0x264E
        "--------", -- 0x264F
        "--------", -- 0x2650
        "--------", -- 0x2651
        "--------", -- 0x2652
        "--------", -- 0x2653
        "--------", -- 0x2654
        "--------", -- 0x2655
        "--------", -- 0x2656
        "--------", -- 0x2657
        "--------", -- 0x2658
        "--------", -- 0x2659
        "--------", -- 0x265A
        "--------", -- 0x265B
        "--------", -- 0x265C
        "--------", -- 0x265D
        "--------", -- 0x265E
        "--------", -- 0x265F
        "--------", -- 0x2660
        "--------", -- 0x2661
        "--------", -- 0x2662
        "--------", -- 0x2663
        "--------", -- 0x2664
        "--------", -- 0x2665
        "--------", -- 0x2666
        "--------", -- 0x2667
        "--------", -- 0x2668
        "--------", -- 0x2669
        "--------", -- 0x266A
        "--------", -- 0x266B
        "--------", -- 0x266C
        "--------", -- 0x266D
        "--------", -- 0x266E
        "--------", -- 0x266F
        "--------", -- 0x2670
        "--------", -- 0x2671
        "--------", -- 0x2672
        "--------", -- 0x2673
        "--------", -- 0x2674
        "--------", -- 0x2675
        "--------", -- 0x2676
        "--------", -- 0x2677
        "--------", -- 0x2678
        "--------", -- 0x2679
        "--------", -- 0x267A
        "--------", -- 0x267B
        "--------", -- 0x267C
        "--------", -- 0x267D
        "--------", -- 0x267E
        "--------", -- 0x267F
        "--------", -- 0x2680
        "--------", -- 0x2681
        "--------", -- 0x2682
        "--------", -- 0x2683
        "--------", -- 0x2684
        "--------", -- 0x2685
        "--------", -- 0x2686
        "--------", -- 0x2687
        "--------", -- 0x2688
        "--------", -- 0x2689
        "--------", -- 0x268A
        "--------", -- 0x268B
        "--------", -- 0x268C
        "--------", -- 0x268D
        "--------", -- 0x268E
        "--------", -- 0x268F
        "--------", -- 0x2690
        "--------", -- 0x2691
        "--------", -- 0x2692
        "--------", -- 0x2693
        "--------", -- 0x2694
        "--------", -- 0x2695
        "--------", -- 0x2696
        "--------", -- 0x2697
        "--------", -- 0x2698
        "--------", -- 0x2699
        "--------", -- 0x269A
        "--------", -- 0x269B
        "--------", -- 0x269C
        "--------", -- 0x269D
        "--------", -- 0x269E
        "--------", -- 0x269F
        "--------", -- 0x26A0
        "--------", -- 0x26A1
        "--------", -- 0x26A2
        "--------", -- 0x26A3
        "--------", -- 0x26A4
        "--------", -- 0x26A5
        "--------", -- 0x26A6
        "--------", -- 0x26A7
        "--------", -- 0x26A8
        "--------", -- 0x26A9
        "--------", -- 0x26AA
        "--------", -- 0x26AB
        "--------", -- 0x26AC
        "--------", -- 0x26AD
        "--------", -- 0x26AE
        "--------", -- 0x26AF
        "--------", -- 0x26B0
        "--------", -- 0x26B1
        "--------", -- 0x26B2
        "--------", -- 0x26B3
        "--------", -- 0x26B4
        "--------", -- 0x26B5
        "--------", -- 0x26B6
        "--------", -- 0x26B7
        "--------", -- 0x26B8
        "--------", -- 0x26B9
        "--------", -- 0x26BA
        "--------", -- 0x26BB
        "--------", -- 0x26BC
        "--------", -- 0x26BD
        "--------", -- 0x26BE
        "--------", -- 0x26BF
        "--------", -- 0x26C0
        "--------", -- 0x26C1
        "--------", -- 0x26C2
        "--------", -- 0x26C3
        "--------", -- 0x26C4
        "--------", -- 0x26C5
        "--------", -- 0x26C6
        "--------", -- 0x26C7
        "--------", -- 0x26C8
        "--------", -- 0x26C9
        "--------", -- 0x26CA
        "--------", -- 0x26CB
        "--------", -- 0x26CC
        "--------", -- 0x26CD
        "--------", -- 0x26CE
        "--------", -- 0x26CF
        "--------", -- 0x26D0
        "--------", -- 0x26D1
        "--------", -- 0x26D2
        "--------", -- 0x26D3
        "--------", -- 0x26D4
        "--------", -- 0x26D5
        "--------", -- 0x26D6
        "--------", -- 0x26D7
        "--------", -- 0x26D8
        "--------", -- 0x26D9
        "--------", -- 0x26DA
        "--------", -- 0x26DB
        "--------", -- 0x26DC
        "--------", -- 0x26DD
        "--------", -- 0x26DE
        "--------", -- 0x26DF
        "--------", -- 0x26E0
        "--------", -- 0x26E1
        "--------", -- 0x26E2
        "--------", -- 0x26E3
        "--------", -- 0x26E4
        "--------", -- 0x26E5
        "--------", -- 0x26E6
        "--------", -- 0x26E7
        "--------", -- 0x26E8
        "--------", -- 0x26E9
        "--------", -- 0x26EA
        "--------", -- 0x26EB
        "--------", -- 0x26EC
        "--------", -- 0x26ED
        "--------", -- 0x26EE
        "--------", -- 0x26EF
        "--------", -- 0x26F0
        "--------", -- 0x26F1
        "--------", -- 0x26F2
        "--------", -- 0x26F3
        "--------", -- 0x26F4
        "--------", -- 0x26F5
        "--------", -- 0x26F6
        "--------", -- 0x26F7
        "--------", -- 0x26F8
        "--------", -- 0x26F9
        "--------", -- 0x26FA
        "--------", -- 0x26FB
        "--------", -- 0x26FC
        "--------", -- 0x26FD
        "--------", -- 0x26FE
        "--------", -- 0x26FF
        "--------", -- 0x2700
        "--------", -- 0x2701
        "--------", -- 0x2702
        "--------", -- 0x2703
        "--------", -- 0x2704
        "--------", -- 0x2705
        "--------", -- 0x2706
        "--------", -- 0x2707
        "--------", -- 0x2708
        "--------", -- 0x2709
        "--------", -- 0x270A
        "--------", -- 0x270B
        "--------", -- 0x270C
        "--------", -- 0x270D
        "--------", -- 0x270E
        "--------", -- 0x270F
        "--------", -- 0x2710
        "--------", -- 0x2711
        "--------", -- 0x2712
        "--------", -- 0x2713
        "--------", -- 0x2714
        "--------", -- 0x2715
        "--------", -- 0x2716
        "--------", -- 0x2717
        "--------", -- 0x2718
        "--------", -- 0x2719
        "--------", -- 0x271A
        "--------", -- 0x271B
        "--------", -- 0x271C
        "--------", -- 0x271D
        "--------", -- 0x271E
        "--------", -- 0x271F
        "--------", -- 0x2720
        "--------", -- 0x2721
        "--------", -- 0x2722
        "--------", -- 0x2723
        "--------", -- 0x2724
        "--------", -- 0x2725
        "--------", -- 0x2726
        "--------", -- 0x2727
        "--------", -- 0x2728
        "--------", -- 0x2729
        "--------", -- 0x272A
        "--------", -- 0x272B
        "--------", -- 0x272C
        "--------", -- 0x272D
        "--------", -- 0x272E
        "--------", -- 0x272F
        "--------", -- 0x2730
        "--------", -- 0x2731
        "--------", -- 0x2732
        "--------", -- 0x2733
        "--------", -- 0x2734
        "--------", -- 0x2735
        "--------", -- 0x2736
        "--------", -- 0x2737
        "--------", -- 0x2738
        "--------", -- 0x2739
        "--------", -- 0x273A
        "--------", -- 0x273B
        "--------", -- 0x273C
        "--------", -- 0x273D
        "--------", -- 0x273E
        "--------", -- 0x273F
        "--------", -- 0x2740
        "--------", -- 0x2741
        "--------", -- 0x2742
        "--------", -- 0x2743
        "--------", -- 0x2744
        "--------", -- 0x2745
        "--------", -- 0x2746
        "--------", -- 0x2747
        "--------", -- 0x2748
        "--------", -- 0x2749
        "--------", -- 0x274A
        "--------", -- 0x274B
        "--------", -- 0x274C
        "--------", -- 0x274D
        "--------", -- 0x274E
        "--------", -- 0x274F
        "--------", -- 0x2750
        "--------", -- 0x2751
        "--------", -- 0x2752
        "--------", -- 0x2753
        "--------", -- 0x2754
        "--------", -- 0x2755
        "--------", -- 0x2756
        "--------", -- 0x2757
        "--------", -- 0x2758
        "--------", -- 0x2759
        "--------", -- 0x275A
        "--------", -- 0x275B
        "--------", -- 0x275C
        "--------", -- 0x275D
        "--------", -- 0x275E
        "--------", -- 0x275F
        "--------", -- 0x2760
        "--------", -- 0x2761
        "--------", -- 0x2762
        "--------", -- 0x2763
        "--------", -- 0x2764
        "--------", -- 0x2765
        "--------", -- 0x2766
        "--------", -- 0x2767
        "--------", -- 0x2768
        "--------", -- 0x2769
        "--------", -- 0x276A
        "--------", -- 0x276B
        "--------", -- 0x276C
        "--------", -- 0x276D
        "--------", -- 0x276E
        "--------", -- 0x276F
        "--------", -- 0x2770
        "--------", -- 0x2771
        "--------", -- 0x2772
        "--------", -- 0x2773
        "--------", -- 0x2774
        "--------", -- 0x2775
        "--------", -- 0x2776
        "--------", -- 0x2777
        "--------", -- 0x2778
        "--------", -- 0x2779
        "--------", -- 0x277A
        "--------", -- 0x277B
        "--------", -- 0x277C
        "--------", -- 0x277D
        "--------", -- 0x277E
        "--------", -- 0x277F
        "--------", -- 0x2780
        "--------", -- 0x2781
        "--------", -- 0x2782
        "--------", -- 0x2783
        "--------", -- 0x2784
        "--------", -- 0x2785
        "--------", -- 0x2786
        "--------", -- 0x2787
        "--------", -- 0x2788
        "--------", -- 0x2789
        "--------", -- 0x278A
        "--------", -- 0x278B
        "--------", -- 0x278C
        "--------", -- 0x278D
        "--------", -- 0x278E
        "--------", -- 0x278F
        "--------", -- 0x2790
        "--------", -- 0x2791
        "--------", -- 0x2792
        "--------", -- 0x2793
        "--------", -- 0x2794
        "--------", -- 0x2795
        "--------", -- 0x2796
        "--------", -- 0x2797
        "--------", -- 0x2798
        "--------", -- 0x2799
        "--------", -- 0x279A
        "--------", -- 0x279B
        "--------", -- 0x279C
        "--------", -- 0x279D
        "--------", -- 0x279E
        "--------", -- 0x279F
        "--------", -- 0x27A0
        "--------", -- 0x27A1
        "--------", -- 0x27A2
        "--------", -- 0x27A3
        "--------", -- 0x27A4
        "--------", -- 0x27A5
        "--------", -- 0x27A6
        "--------", -- 0x27A7
        "--------", -- 0x27A8
        "--------", -- 0x27A9
        "--------", -- 0x27AA
        "--------", -- 0x27AB
        "--------", -- 0x27AC
        "--------", -- 0x27AD
        "--------", -- 0x27AE
        "--------", -- 0x27AF
        "--------", -- 0x27B0
        "--------", -- 0x27B1
        "--------", -- 0x27B2
        "--------", -- 0x27B3
        "--------", -- 0x27B4
        "--------", -- 0x27B5
        "--------", -- 0x27B6
        "--------", -- 0x27B7
        "--------", -- 0x27B8
        "--------", -- 0x27B9
        "--------", -- 0x27BA
        "--------", -- 0x27BB
        "--------", -- 0x27BC
        "--------", -- 0x27BD
        "--------", -- 0x27BE
        "--------", -- 0x27BF
        "--------", -- 0x27C0
        "--------", -- 0x27C1
        "--------", -- 0x27C2
        "--------", -- 0x27C3
        "--------", -- 0x27C4
        "--------", -- 0x27C5
        "--------", -- 0x27C6
        "--------", -- 0x27C7
        "--------", -- 0x27C8
        "--------", -- 0x27C9
        "--------", -- 0x27CA
        "--------", -- 0x27CB
        "--------", -- 0x27CC
        "--------", -- 0x27CD
        "--------", -- 0x27CE
        "--------", -- 0x27CF
        "--------", -- 0x27D0
        "--------", -- 0x27D1
        "--------", -- 0x27D2
        "--------", -- 0x27D3
        "--------", -- 0x27D4
        "--------", -- 0x27D5
        "--------", -- 0x27D6
        "--------", -- 0x27D7
        "--------", -- 0x27D8
        "--------", -- 0x27D9
        "--------", -- 0x27DA
        "--------", -- 0x27DB
        "--------", -- 0x27DC
        "--------", -- 0x27DD
        "--------", -- 0x27DE
        "--------", -- 0x27DF
        "--------", -- 0x27E0
        "--------", -- 0x27E1
        "--------", -- 0x27E2
        "--------", -- 0x27E3
        "--------", -- 0x27E4
        "--------", -- 0x27E5
        "--------", -- 0x27E6
        "--------", -- 0x27E7
        "--------", -- 0x27E8
        "--------", -- 0x27E9
        "--------", -- 0x27EA
        "--------", -- 0x27EB
        "--------", -- 0x27EC
        "--------", -- 0x27ED
        "--------", -- 0x27EE
        "--------", -- 0x27EF
        "--------", -- 0x27F0
        "--------", -- 0x27F1
        "--------", -- 0x27F2
        "--------", -- 0x27F3
        "--------", -- 0x27F4
        "--------", -- 0x27F5
        "--------", -- 0x27F6
        "--------", -- 0x27F7
        "--------", -- 0x27F8
        "--------", -- 0x27F9
        "--------", -- 0x27FA
        "--------", -- 0x27FB
        "--------", -- 0x27FC
        "--------", -- 0x27FD
        "--------", -- 0x27FE
        "--------", -- 0x27FF
        "--------", -- 0x2800
        "--------", -- 0x2801
        "--------", -- 0x2802
        "--------", -- 0x2803
        "--------", -- 0x2804
        "--------", -- 0x2805
        "--------", -- 0x2806
        "--------", -- 0x2807
        "--------", -- 0x2808
        "--------", -- 0x2809
        "--------", -- 0x280A
        "--------", -- 0x280B
        "--------", -- 0x280C
        "--------", -- 0x280D
        "--------", -- 0x280E
        "--------", -- 0x280F
        "--------", -- 0x2810
        "--------", -- 0x2811
        "--------", -- 0x2812
        "--------", -- 0x2813
        "--------", -- 0x2814
        "--------", -- 0x2815
        "--------", -- 0x2816
        "--------", -- 0x2817
        "--------", -- 0x2818
        "--------", -- 0x2819
        "--------", -- 0x281A
        "--------", -- 0x281B
        "--------", -- 0x281C
        "--------", -- 0x281D
        "--------", -- 0x281E
        "--------", -- 0x281F
        "--------", -- 0x2820
        "--------", -- 0x2821
        "--------", -- 0x2822
        "--------", -- 0x2823
        "--------", -- 0x2824
        "--------", -- 0x2825
        "--------", -- 0x2826
        "--------", -- 0x2827
        "--------", -- 0x2828
        "--------", -- 0x2829
        "--------", -- 0x282A
        "--------", -- 0x282B
        "--------", -- 0x282C
        "--------", -- 0x282D
        "--------", -- 0x282E
        "--------", -- 0x282F
        "--------", -- 0x2830
        "--------", -- 0x2831
        "--------", -- 0x2832
        "--------", -- 0x2833
        "--------", -- 0x2834
        "--------", -- 0x2835
        "--------", -- 0x2836
        "--------", -- 0x2837
        "--------", -- 0x2838
        "--------", -- 0x2839
        "--------", -- 0x283A
        "--------", -- 0x283B
        "--------", -- 0x283C
        "--------", -- 0x283D
        "--------", -- 0x283E
        "--------", -- 0x283F
        "--------", -- 0x2840
        "--------", -- 0x2841
        "--------", -- 0x2842
        "--------", -- 0x2843
        "--------", -- 0x2844
        "--------", -- 0x2845
        "--------", -- 0x2846
        "--------", -- 0x2847
        "--------", -- 0x2848
        "--------", -- 0x2849
        "--------", -- 0x284A
        "--------", -- 0x284B
        "--------", -- 0x284C
        "--------", -- 0x284D
        "--------", -- 0x284E
        "--------", -- 0x284F
        "--------", -- 0x2850
        "--------", -- 0x2851
        "--------", -- 0x2852
        "--------", -- 0x2853
        "--------", -- 0x2854
        "--------", -- 0x2855
        "--------", -- 0x2856
        "--------", -- 0x2857
        "--------", -- 0x2858
        "--------", -- 0x2859
        "--------", -- 0x285A
        "--------", -- 0x285B
        "--------", -- 0x285C
        "--------", -- 0x285D
        "--------", -- 0x285E
        "--------", -- 0x285F
        "--------", -- 0x2860
        "--------", -- 0x2861
        "--------", -- 0x2862
        "--------", -- 0x2863
        "--------", -- 0x2864
        "--------", -- 0x2865
        "--------", -- 0x2866
        "--------", -- 0x2867
        "--------", -- 0x2868
        "--------", -- 0x2869
        "--------", -- 0x286A
        "--------", -- 0x286B
        "--------", -- 0x286C
        "--------", -- 0x286D
        "--------", -- 0x286E
        "--------", -- 0x286F
        "--------", -- 0x2870
        "--------", -- 0x2871
        "--------", -- 0x2872
        "--------", -- 0x2873
        "--------", -- 0x2874
        "--------", -- 0x2875
        "--------", -- 0x2876
        "--------", -- 0x2877
        "--------", -- 0x2878
        "--------", -- 0x2879
        "--------", -- 0x287A
        "--------", -- 0x287B
        "--------", -- 0x287C
        "--------", -- 0x287D
        "--------", -- 0x287E
        "--------", -- 0x287F
        "--------", -- 0x2880
        "--------", -- 0x2881
        "--------", -- 0x2882
        "--------", -- 0x2883
        "--------", -- 0x2884
        "--------", -- 0x2885
        "--------", -- 0x2886
        "--------", -- 0x2887
        "--------", -- 0x2888
        "--------", -- 0x2889
        "--------", -- 0x288A
        "--------", -- 0x288B
        "--------", -- 0x288C
        "--------", -- 0x288D
        "--------", -- 0x288E
        "--------", -- 0x288F
        "--------", -- 0x2890
        "--------", -- 0x2891
        "--------", -- 0x2892
        "--------", -- 0x2893
        "--------", -- 0x2894
        "--------", -- 0x2895
        "--------", -- 0x2896
        "--------", -- 0x2897
        "--------", -- 0x2898
        "--------", -- 0x2899
        "--------", -- 0x289A
        "--------", -- 0x289B
        "--------", -- 0x289C
        "--------", -- 0x289D
        "--------", -- 0x289E
        "--------", -- 0x289F
        "--------", -- 0x28A0
        "--------", -- 0x28A1
        "--------", -- 0x28A2
        "--------", -- 0x28A3
        "--------", -- 0x28A4
        "--------", -- 0x28A5
        "--------", -- 0x28A6
        "--------", -- 0x28A7
        "--------", -- 0x28A8
        "--------", -- 0x28A9
        "--------", -- 0x28AA
        "--------", -- 0x28AB
        "--------", -- 0x28AC
        "--------", -- 0x28AD
        "--------", -- 0x28AE
        "--------", -- 0x28AF
        "--------", -- 0x28B0
        "--------", -- 0x28B1
        "--------", -- 0x28B2
        "--------", -- 0x28B3
        "--------", -- 0x28B4
        "--------", -- 0x28B5
        "--------", -- 0x28B6
        "--------", -- 0x28B7
        "--------", -- 0x28B8
        "--------", -- 0x28B9
        "--------", -- 0x28BA
        "--------", -- 0x28BB
        "--------", -- 0x28BC
        "--------", -- 0x28BD
        "--------", -- 0x28BE
        "--------", -- 0x28BF
        "--------", -- 0x28C0
        "--------", -- 0x28C1
        "--------", -- 0x28C2
        "--------", -- 0x28C3
        "--------", -- 0x28C4
        "--------", -- 0x28C5
        "--------", -- 0x28C6
        "--------", -- 0x28C7
        "--------", -- 0x28C8
        "--------", -- 0x28C9
        "--------", -- 0x28CA
        "--------", -- 0x28CB
        "--------", -- 0x28CC
        "--------", -- 0x28CD
        "--------", -- 0x28CE
        "--------", -- 0x28CF
        "--------", -- 0x28D0
        "--------", -- 0x28D1
        "--------", -- 0x28D2
        "--------", -- 0x28D3
        "--------", -- 0x28D4
        "--------", -- 0x28D5
        "--------", -- 0x28D6
        "--------", -- 0x28D7
        "--------", -- 0x28D8
        "--------", -- 0x28D9
        "--------", -- 0x28DA
        "--------", -- 0x28DB
        "--------", -- 0x28DC
        "--------", -- 0x28DD
        "--------", -- 0x28DE
        "--------", -- 0x28DF
        "--------", -- 0x28E0
        "--------", -- 0x28E1
        "--------", -- 0x28E2
        "--------", -- 0x28E3
        "--------", -- 0x28E4
        "--------", -- 0x28E5
        "--------", -- 0x28E6
        "--------", -- 0x28E7
        "--------", -- 0x28E8
        "--------", -- 0x28E9
        "--------", -- 0x28EA
        "--------", -- 0x28EB
        "--------", -- 0x28EC
        "--------", -- 0x28ED
        "--------", -- 0x28EE
        "--------", -- 0x28EF
        "--------", -- 0x28F0
        "--------", -- 0x28F1
        "--------", -- 0x28F2
        "--------", -- 0x28F3
        "--------", -- 0x28F4
        "--------", -- 0x28F5
        "--------", -- 0x28F6
        "--------", -- 0x28F7
        "--------", -- 0x28F8
        "--------", -- 0x28F9
        "--------", -- 0x28FA
        "--------", -- 0x28FB
        "--------", -- 0x28FC
        "--------", -- 0x28FD
        "--------", -- 0x28FE
        "--------", -- 0x28FF
        "--------", -- 0x2900
        "--------", -- 0x2901
        "--------", -- 0x2902
        "--------", -- 0x2903
        "--------", -- 0x2904
        "--------", -- 0x2905
        "--------", -- 0x2906
        "--------", -- 0x2907
        "--------", -- 0x2908
        "--------", -- 0x2909
        "--------", -- 0x290A
        "--------", -- 0x290B
        "--------", -- 0x290C
        "--------", -- 0x290D
        "--------", -- 0x290E
        "--------", -- 0x290F
        "--------", -- 0x2910
        "--------", -- 0x2911
        "--------", -- 0x2912
        "--------", -- 0x2913
        "--------", -- 0x2914
        "--------", -- 0x2915
        "--------", -- 0x2916
        "--------", -- 0x2917
        "--------", -- 0x2918
        "--------", -- 0x2919
        "--------", -- 0x291A
        "--------", -- 0x291B
        "--------", -- 0x291C
        "--------", -- 0x291D
        "--------", -- 0x291E
        "--------", -- 0x291F
        "--------", -- 0x2920
        "--------", -- 0x2921
        "--------", -- 0x2922
        "--------", -- 0x2923
        "--------", -- 0x2924
        "--------", -- 0x2925
        "--------", -- 0x2926
        "--------", -- 0x2927
        "--------", -- 0x2928
        "--------", -- 0x2929
        "--------", -- 0x292A
        "--------", -- 0x292B
        "--------", -- 0x292C
        "--------", -- 0x292D
        "--------", -- 0x292E
        "--------", -- 0x292F
        "--------", -- 0x2930
        "--------", -- 0x2931
        "--------", -- 0x2932
        "--------", -- 0x2933
        "--------", -- 0x2934
        "--------", -- 0x2935
        "--------", -- 0x2936
        "--------", -- 0x2937
        "--------", -- 0x2938
        "--------", -- 0x2939
        "--------", -- 0x293A
        "--------", -- 0x293B
        "--------", -- 0x293C
        "--------", -- 0x293D
        "--------", -- 0x293E
        "--------", -- 0x293F
        "--------", -- 0x2940
        "--------", -- 0x2941
        "--------", -- 0x2942
        "--------", -- 0x2943
        "--------", -- 0x2944
        "--------", -- 0x2945
        "--------", -- 0x2946
        "--------", -- 0x2947
        "--------", -- 0x2948
        "--------", -- 0x2949
        "--------", -- 0x294A
        "--------", -- 0x294B
        "--------", -- 0x294C
        "--------", -- 0x294D
        "--------", -- 0x294E
        "--------", -- 0x294F
        "--------", -- 0x2950
        "--------", -- 0x2951
        "--------", -- 0x2952
        "--------", -- 0x2953
        "--------", -- 0x2954
        "--------", -- 0x2955
        "--------", -- 0x2956
        "--------", -- 0x2957
        "--------", -- 0x2958
        "--------", -- 0x2959
        "--------", -- 0x295A
        "--------", -- 0x295B
        "--------", -- 0x295C
        "--------", -- 0x295D
        "--------", -- 0x295E
        "--------", -- 0x295F
        "--------", -- 0x2960
        "--------", -- 0x2961
        "--------", -- 0x2962
        "--------", -- 0x2963
        "--------", -- 0x2964
        "--------", -- 0x2965
        "--------", -- 0x2966
        "--------", -- 0x2967
        "--------", -- 0x2968
        "--------", -- 0x2969
        "--------", -- 0x296A
        "--------", -- 0x296B
        "--------", -- 0x296C
        "--------", -- 0x296D
        "--------", -- 0x296E
        "--------", -- 0x296F
        "--------", -- 0x2970
        "--------", -- 0x2971
        "--------", -- 0x2972
        "--------", -- 0x2973
        "--------", -- 0x2974
        "--------", -- 0x2975
        "--------", -- 0x2976
        "--------", -- 0x2977
        "--------", -- 0x2978
        "--------", -- 0x2979
        "--------", -- 0x297A
        "--------", -- 0x297B
        "--------", -- 0x297C
        "--------", -- 0x297D
        "--------", -- 0x297E
        "--------", -- 0x297F
        "--------", -- 0x2980
        "--------", -- 0x2981
        "--------", -- 0x2982
        "--------", -- 0x2983
        "--------", -- 0x2984
        "--------", -- 0x2985
        "--------", -- 0x2986
        "--------", -- 0x2987
        "--------", -- 0x2988
        "--------", -- 0x2989
        "--------", -- 0x298A
        "--------", -- 0x298B
        "--------", -- 0x298C
        "--------", -- 0x298D
        "--------", -- 0x298E
        "--------", -- 0x298F
        "--------", -- 0x2990
        "--------", -- 0x2991
        "--------", -- 0x2992
        "--------", -- 0x2993
        "--------", -- 0x2994
        "--------", -- 0x2995
        "--------", -- 0x2996
        "--------", -- 0x2997
        "--------", -- 0x2998
        "--------", -- 0x2999
        "--------", -- 0x299A
        "--------", -- 0x299B
        "--------", -- 0x299C
        "--------", -- 0x299D
        "--------", -- 0x299E
        "--------", -- 0x299F
        "--------", -- 0x29A0
        "--------", -- 0x29A1
        "--------", -- 0x29A2
        "--------", -- 0x29A3
        "--------", -- 0x29A4
        "--------", -- 0x29A5
        "--------", -- 0x29A6
        "--------", -- 0x29A7
        "--------", -- 0x29A8
        "--------", -- 0x29A9
        "--------", -- 0x29AA
        "--------", -- 0x29AB
        "--------", -- 0x29AC
        "--------", -- 0x29AD
        "--------", -- 0x29AE
        "--------", -- 0x29AF
        "--------", -- 0x29B0
        "--------", -- 0x29B1
        "--------", -- 0x29B2
        "--------", -- 0x29B3
        "--------", -- 0x29B4
        "--------", -- 0x29B5
        "--------", -- 0x29B6
        "--------", -- 0x29B7
        "--------", -- 0x29B8
        "--------", -- 0x29B9
        "--------", -- 0x29BA
        "--------", -- 0x29BB
        "--------", -- 0x29BC
        "--------", -- 0x29BD
        "--------", -- 0x29BE
        "--------", -- 0x29BF
        "--------", -- 0x29C0
        "--------", -- 0x29C1
        "--------", -- 0x29C2
        "--------", -- 0x29C3
        "--------", -- 0x29C4
        "--------", -- 0x29C5
        "--------", -- 0x29C6
        "--------", -- 0x29C7
        "--------", -- 0x29C8
        "--------", -- 0x29C9
        "--------", -- 0x29CA
        "--------", -- 0x29CB
        "--------", -- 0x29CC
        "--------", -- 0x29CD
        "--------", -- 0x29CE
        "--------", -- 0x29CF
        "--------", -- 0x29D0
        "--------", -- 0x29D1
        "--------", -- 0x29D2
        "--------", -- 0x29D3
        "--------", -- 0x29D4
        "--------", -- 0x29D5
        "--------", -- 0x29D6
        "--------", -- 0x29D7
        "--------", -- 0x29D8
        "--------", -- 0x29D9
        "--------", -- 0x29DA
        "--------", -- 0x29DB
        "--------", -- 0x29DC
        "--------", -- 0x29DD
        "--------", -- 0x29DE
        "--------", -- 0x29DF
        "--------", -- 0x29E0
        "--------", -- 0x29E1
        "--------", -- 0x29E2
        "--------", -- 0x29E3
        "--------", -- 0x29E4
        "--------", -- 0x29E5
        "--------", -- 0x29E6
        "--------", -- 0x29E7
        "--------", -- 0x29E8
        "--------", -- 0x29E9
        "--------", -- 0x29EA
        "--------", -- 0x29EB
        "--------", -- 0x29EC
        "--------", -- 0x29ED
        "--------", -- 0x29EE
        "--------", -- 0x29EF
        "--------", -- 0x29F0
        "--------", -- 0x29F1
        "--------", -- 0x29F2
        "--------", -- 0x29F3
        "--------", -- 0x29F4
        "--------", -- 0x29F5
        "--------", -- 0x29F6
        "--------", -- 0x29F7
        "--------", -- 0x29F8
        "--------", -- 0x29F9
        "--------", -- 0x29FA
        "--------", -- 0x29FB
        "--------", -- 0x29FC
        "--------", -- 0x29FD
        "--------", -- 0x29FE
        "--------", -- 0x29FF
        "--------", -- 0x2A00
        "--------", -- 0x2A01
        "--------", -- 0x2A02
        "--------", -- 0x2A03
        "--------", -- 0x2A04
        "--------", -- 0x2A05
        "--------", -- 0x2A06
        "--------", -- 0x2A07
        "--------", -- 0x2A08
        "--------", -- 0x2A09
        "--------", -- 0x2A0A
        "--------", -- 0x2A0B
        "--------", -- 0x2A0C
        "--------", -- 0x2A0D
        "--------", -- 0x2A0E
        "--------", -- 0x2A0F
        "--------", -- 0x2A10
        "--------", -- 0x2A11
        "--------", -- 0x2A12
        "--------", -- 0x2A13
        "--------", -- 0x2A14
        "--------", -- 0x2A15
        "--------", -- 0x2A16
        "--------", -- 0x2A17
        "--------", -- 0x2A18
        "--------", -- 0x2A19
        "--------", -- 0x2A1A
        "--------", -- 0x2A1B
        "--------", -- 0x2A1C
        "--------", -- 0x2A1D
        "--------", -- 0x2A1E
        "--------", -- 0x2A1F
        "--------", -- 0x2A20
        "--------", -- 0x2A21
        "--------", -- 0x2A22
        "--------", -- 0x2A23
        "--------", -- 0x2A24
        "--------", -- 0x2A25
        "--------", -- 0x2A26
        "--------", -- 0x2A27
        "--------", -- 0x2A28
        "--------", -- 0x2A29
        "--------", -- 0x2A2A
        "--------", -- 0x2A2B
        "--------", -- 0x2A2C
        "--------", -- 0x2A2D
        "--------", -- 0x2A2E
        "--------", -- 0x2A2F
        "--------", -- 0x2A30
        "--------", -- 0x2A31
        "--------", -- 0x2A32
        "--------", -- 0x2A33
        "--------", -- 0x2A34
        "--------", -- 0x2A35
        "--------", -- 0x2A36
        "--------", -- 0x2A37
        "--------", -- 0x2A38
        "--------", -- 0x2A39
        "--------", -- 0x2A3A
        "--------", -- 0x2A3B
        "--------", -- 0x2A3C
        "--------", -- 0x2A3D
        "--------", -- 0x2A3E
        "--------", -- 0x2A3F
        "--------", -- 0x2A40
        "--------", -- 0x2A41
        "--------", -- 0x2A42
        "--------", -- 0x2A43
        "--------", -- 0x2A44
        "--------", -- 0x2A45
        "--------", -- 0x2A46
        "--------", -- 0x2A47
        "--------", -- 0x2A48
        "--------", -- 0x2A49
        "--------", -- 0x2A4A
        "--------", -- 0x2A4B
        "--------", -- 0x2A4C
        "--------", -- 0x2A4D
        "--------", -- 0x2A4E
        "--------", -- 0x2A4F
        "--------", -- 0x2A50
        "--------", -- 0x2A51
        "--------", -- 0x2A52
        "--------", -- 0x2A53
        "--------", -- 0x2A54
        "--------", -- 0x2A55
        "--------", -- 0x2A56
        "--------", -- 0x2A57
        "--------", -- 0x2A58
        "--------", -- 0x2A59
        "--------", -- 0x2A5A
        "--------", -- 0x2A5B
        "--------", -- 0x2A5C
        "--------", -- 0x2A5D
        "--------", -- 0x2A5E
        "--------", -- 0x2A5F
        "--------", -- 0x2A60
        "--------", -- 0x2A61
        "--------", -- 0x2A62
        "--------", -- 0x2A63
        "--------", -- 0x2A64
        "--------", -- 0x2A65
        "--------", -- 0x2A66
        "--------", -- 0x2A67
        "--------", -- 0x2A68
        "--------", -- 0x2A69
        "--------", -- 0x2A6A
        "--------", -- 0x2A6B
        "--------", -- 0x2A6C
        "--------", -- 0x2A6D
        "--------", -- 0x2A6E
        "--------", -- 0x2A6F
        "--------", -- 0x2A70
        "--------", -- 0x2A71
        "--------", -- 0x2A72
        "--------", -- 0x2A73
        "--------", -- 0x2A74
        "--------", -- 0x2A75
        "--------", -- 0x2A76
        "--------", -- 0x2A77
        "--------", -- 0x2A78
        "--------", -- 0x2A79
        "--------", -- 0x2A7A
        "--------", -- 0x2A7B
        "--------", -- 0x2A7C
        "--------", -- 0x2A7D
        "--------", -- 0x2A7E
        "--------", -- 0x2A7F
        "--------", -- 0x2A80
        "--------", -- 0x2A81
        "--------", -- 0x2A82
        "--------", -- 0x2A83
        "--------", -- 0x2A84
        "--------", -- 0x2A85
        "--------", -- 0x2A86
        "--------", -- 0x2A87
        "--------", -- 0x2A88
        "--------", -- 0x2A89
        "--------", -- 0x2A8A
        "--------", -- 0x2A8B
        "--------", -- 0x2A8C
        "--------", -- 0x2A8D
        "--------", -- 0x2A8E
        "--------", -- 0x2A8F
        "--------", -- 0x2A90
        "--------", -- 0x2A91
        "--------", -- 0x2A92
        "--------", -- 0x2A93
        "--------", -- 0x2A94
        "--------", -- 0x2A95
        "--------", -- 0x2A96
        "--------", -- 0x2A97
        "--------", -- 0x2A98
        "--------", -- 0x2A99
        "--------", -- 0x2A9A
        "--------", -- 0x2A9B
        "--------", -- 0x2A9C
        "--------", -- 0x2A9D
        "--------", -- 0x2A9E
        "--------", -- 0x2A9F
        "--------", -- 0x2AA0
        "--------", -- 0x2AA1
        "--------", -- 0x2AA2
        "--------", -- 0x2AA3
        "--------", -- 0x2AA4
        "--------", -- 0x2AA5
        "--------", -- 0x2AA6
        "--------", -- 0x2AA7
        "--------", -- 0x2AA8
        "--------", -- 0x2AA9
        "--------", -- 0x2AAA
        "--------", -- 0x2AAB
        "--------", -- 0x2AAC
        "--------", -- 0x2AAD
        "--------", -- 0x2AAE
        "--------", -- 0x2AAF
        "--------", -- 0x2AB0
        "--------", -- 0x2AB1
        "--------", -- 0x2AB2
        "--------", -- 0x2AB3
        "--------", -- 0x2AB4
        "--------", -- 0x2AB5
        "--------", -- 0x2AB6
        "--------", -- 0x2AB7
        "--------", -- 0x2AB8
        "--------", -- 0x2AB9
        "--------", -- 0x2ABA
        "--------", -- 0x2ABB
        "--------", -- 0x2ABC
        "--------", -- 0x2ABD
        "--------", -- 0x2ABE
        "--------", -- 0x2ABF
        "--------", -- 0x2AC0
        "--------", -- 0x2AC1
        "--------", -- 0x2AC2
        "--------", -- 0x2AC3
        "--------", -- 0x2AC4
        "--------", -- 0x2AC5
        "--------", -- 0x2AC6
        "--------", -- 0x2AC7
        "--------", -- 0x2AC8
        "--------", -- 0x2AC9
        "--------", -- 0x2ACA
        "--------", -- 0x2ACB
        "--------", -- 0x2ACC
        "--------", -- 0x2ACD
        "--------", -- 0x2ACE
        "--------", -- 0x2ACF
        "--------", -- 0x2AD0
        "--------", -- 0x2AD1
        "--------", -- 0x2AD2
        "--------", -- 0x2AD3
        "--------", -- 0x2AD4
        "--------", -- 0x2AD5
        "--------", -- 0x2AD6
        "--------", -- 0x2AD7
        "--------", -- 0x2AD8
        "--------", -- 0x2AD9
        "--------", -- 0x2ADA
        "--------", -- 0x2ADB
        "--------", -- 0x2ADC
        "--------", -- 0x2ADD
        "--------", -- 0x2ADE
        "--------", -- 0x2ADF
        "--------", -- 0x2AE0
        "--------", -- 0x2AE1
        "--------", -- 0x2AE2
        "--------", -- 0x2AE3
        "--------", -- 0x2AE4
        "--------", -- 0x2AE5
        "--------", -- 0x2AE6
        "--------", -- 0x2AE7
        "--------", -- 0x2AE8
        "--------", -- 0x2AE9
        "--------", -- 0x2AEA
        "--------", -- 0x2AEB
        "--------", -- 0x2AEC
        "--------", -- 0x2AED
        "--------", -- 0x2AEE
        "--------", -- 0x2AEF
        "--------", -- 0x2AF0
        "--------", -- 0x2AF1
        "--------", -- 0x2AF2
        "--------", -- 0x2AF3
        "--------", -- 0x2AF4
        "--------", -- 0x2AF5
        "--------", -- 0x2AF6
        "--------", -- 0x2AF7
        "--------", -- 0x2AF8
        "--------", -- 0x2AF9
        "--------", -- 0x2AFA
        "--------", -- 0x2AFB
        "--------", -- 0x2AFC
        "--------", -- 0x2AFD
        "--------", -- 0x2AFE
        "--------", -- 0x2AFF
        "--------", -- 0x2B00
        "--------", -- 0x2B01
        "--------", -- 0x2B02
        "--------", -- 0x2B03
        "--------", -- 0x2B04
        "--------", -- 0x2B05
        "--------", -- 0x2B06
        "--------", -- 0x2B07
        "--------", -- 0x2B08
        "--------", -- 0x2B09
        "--------", -- 0x2B0A
        "--------", -- 0x2B0B
        "--------", -- 0x2B0C
        "--------", -- 0x2B0D
        "--------", -- 0x2B0E
        "--------", -- 0x2B0F
        "--------", -- 0x2B10
        "--------", -- 0x2B11
        "--------", -- 0x2B12
        "--------", -- 0x2B13
        "--------", -- 0x2B14
        "--------", -- 0x2B15
        "--------", -- 0x2B16
        "--------", -- 0x2B17
        "--------", -- 0x2B18
        "--------", -- 0x2B19
        "--------", -- 0x2B1A
        "--------", -- 0x2B1B
        "--------", -- 0x2B1C
        "--------", -- 0x2B1D
        "--------", -- 0x2B1E
        "--------", -- 0x2B1F
        "--------", -- 0x2B20
        "--------", -- 0x2B21
        "--------", -- 0x2B22
        "--------", -- 0x2B23
        "--------", -- 0x2B24
        "--------", -- 0x2B25
        "--------", -- 0x2B26
        "--------", -- 0x2B27
        "--------", -- 0x2B28
        "--------", -- 0x2B29
        "--------", -- 0x2B2A
        "--------", -- 0x2B2B
        "--------", -- 0x2B2C
        "--------", -- 0x2B2D
        "--------", -- 0x2B2E
        "--------", -- 0x2B2F
        "--------", -- 0x2B30
        "--------", -- 0x2B31
        "--------", -- 0x2B32
        "--------", -- 0x2B33
        "--------", -- 0x2B34
        "--------", -- 0x2B35
        "--------", -- 0x2B36
        "--------", -- 0x2B37
        "--------", -- 0x2B38
        "--------", -- 0x2B39
        "--------", -- 0x2B3A
        "--------", -- 0x2B3B
        "--------", -- 0x2B3C
        "--------", -- 0x2B3D
        "--------", -- 0x2B3E
        "--------", -- 0x2B3F
        "--------", -- 0x2B40
        "--------", -- 0x2B41
        "--------", -- 0x2B42
        "--------", -- 0x2B43
        "--------", -- 0x2B44
        "--------", -- 0x2B45
        "--------", -- 0x2B46
        "--------", -- 0x2B47
        "--------", -- 0x2B48
        "--------", -- 0x2B49
        "--------", -- 0x2B4A
        "--------", -- 0x2B4B
        "--------", -- 0x2B4C
        "--------", -- 0x2B4D
        "--------", -- 0x2B4E
        "--------", -- 0x2B4F
        "--------", -- 0x2B50
        "--------", -- 0x2B51
        "--------", -- 0x2B52
        "--------", -- 0x2B53
        "--------", -- 0x2B54
        "--------", -- 0x2B55
        "--------", -- 0x2B56
        "--------", -- 0x2B57
        "--------", -- 0x2B58
        "--------", -- 0x2B59
        "--------", -- 0x2B5A
        "--------", -- 0x2B5B
        "--------", -- 0x2B5C
        "--------", -- 0x2B5D
        "--------", -- 0x2B5E
        "--------", -- 0x2B5F
        "--------", -- 0x2B60
        "--------", -- 0x2B61
        "--------", -- 0x2B62
        "--------", -- 0x2B63
        "--------", -- 0x2B64
        "--------", -- 0x2B65
        "--------", -- 0x2B66
        "--------", -- 0x2B67
        "--------", -- 0x2B68
        "--------", -- 0x2B69
        "--------", -- 0x2B6A
        "--------", -- 0x2B6B
        "--------", -- 0x2B6C
        "--------", -- 0x2B6D
        "--------", -- 0x2B6E
        "--------", -- 0x2B6F
        "--------", -- 0x2B70
        "--------", -- 0x2B71
        "--------", -- 0x2B72
        "--------", -- 0x2B73
        "--------", -- 0x2B74
        "--------", -- 0x2B75
        "--------", -- 0x2B76
        "--------", -- 0x2B77
        "--------", -- 0x2B78
        "--------", -- 0x2B79
        "--------", -- 0x2B7A
        "--------", -- 0x2B7B
        "--------", -- 0x2B7C
        "--------", -- 0x2B7D
        "--------", -- 0x2B7E
        "--------", -- 0x2B7F
        "--------", -- 0x2B80
        "--------", -- 0x2B81
        "--------", -- 0x2B82
        "--------", -- 0x2B83
        "--------", -- 0x2B84
        "--------", -- 0x2B85
        "--------", -- 0x2B86
        "--------", -- 0x2B87
        "--------", -- 0x2B88
        "--------", -- 0x2B89
        "--------", -- 0x2B8A
        "--------", -- 0x2B8B
        "--------", -- 0x2B8C
        "--------", -- 0x2B8D
        "--------", -- 0x2B8E
        "--------", -- 0x2B8F
        "--------", -- 0x2B90
        "--------", -- 0x2B91
        "--------", -- 0x2B92
        "--------", -- 0x2B93
        "--------", -- 0x2B94
        "--------", -- 0x2B95
        "--------", -- 0x2B96
        "--------", -- 0x2B97
        "--------", -- 0x2B98
        "--------", -- 0x2B99
        "--------", -- 0x2B9A
        "--------", -- 0x2B9B
        "--------", -- 0x2B9C
        "--------", -- 0x2B9D
        "--------", -- 0x2B9E
        "--------", -- 0x2B9F
        "--------", -- 0x2BA0
        "--------", -- 0x2BA1
        "--------", -- 0x2BA2
        "--------", -- 0x2BA3
        "--------", -- 0x2BA4
        "--------", -- 0x2BA5
        "--------", -- 0x2BA6
        "--------", -- 0x2BA7
        "--------", -- 0x2BA8
        "--------", -- 0x2BA9
        "--------", -- 0x2BAA
        "--------", -- 0x2BAB
        "--------", -- 0x2BAC
        "--------", -- 0x2BAD
        "--------", -- 0x2BAE
        "--------", -- 0x2BAF
        "--------", -- 0x2BB0
        "--------", -- 0x2BB1
        "--------", -- 0x2BB2
        "--------", -- 0x2BB3
        "--------", -- 0x2BB4
        "--------", -- 0x2BB5
        "--------", -- 0x2BB6
        "--------", -- 0x2BB7
        "--------", -- 0x2BB8
        "--------", -- 0x2BB9
        "--------", -- 0x2BBA
        "--------", -- 0x2BBB
        "--------", -- 0x2BBC
        "--------", -- 0x2BBD
        "--------", -- 0x2BBE
        "--------", -- 0x2BBF
        "--------", -- 0x2BC0
        "--------", -- 0x2BC1
        "--------", -- 0x2BC2
        "--------", -- 0x2BC3
        "--------", -- 0x2BC4
        "--------", -- 0x2BC5
        "--------", -- 0x2BC6
        "--------", -- 0x2BC7
        "--------", -- 0x2BC8
        "--------", -- 0x2BC9
        "--------", -- 0x2BCA
        "--------", -- 0x2BCB
        "--------", -- 0x2BCC
        "--------", -- 0x2BCD
        "--------", -- 0x2BCE
        "--------", -- 0x2BCF
        "--------", -- 0x2BD0
        "--------", -- 0x2BD1
        "--------", -- 0x2BD2
        "--------", -- 0x2BD3
        "--------", -- 0x2BD4
        "--------", -- 0x2BD5
        "--------", -- 0x2BD6
        "--------", -- 0x2BD7
        "--------", -- 0x2BD8
        "--------", -- 0x2BD9
        "--------", -- 0x2BDA
        "--------", -- 0x2BDB
        "--------", -- 0x2BDC
        "--------", -- 0x2BDD
        "--------", -- 0x2BDE
        "--------", -- 0x2BDF
        "--------", -- 0x2BE0
        "--------", -- 0x2BE1
        "--------", -- 0x2BE2
        "--------", -- 0x2BE3
        "--------", -- 0x2BE4
        "--------", -- 0x2BE5
        "--------", -- 0x2BE6
        "--------", -- 0x2BE7
        "--------", -- 0x2BE8
        "--------", -- 0x2BE9
        "--------", -- 0x2BEA
        "--------", -- 0x2BEB
        "--------", -- 0x2BEC
        "--------", -- 0x2BED
        "--------", -- 0x2BEE
        "--------", -- 0x2BEF
        "--------", -- 0x2BF0
        "--------", -- 0x2BF1
        "--------", -- 0x2BF2
        "--------", -- 0x2BF3
        "--------", -- 0x2BF4
        "--------", -- 0x2BF5
        "--------", -- 0x2BF6
        "--------", -- 0x2BF7
        "--------", -- 0x2BF8
        "--------", -- 0x2BF9
        "--------", -- 0x2BFA
        "--------", -- 0x2BFB
        "--------", -- 0x2BFC
        "--------", -- 0x2BFD
        "--------", -- 0x2BFE
        "--------", -- 0x2BFF
        "--------", -- 0x2C00
        "--------", -- 0x2C01
        "--------", -- 0x2C02
        "--------", -- 0x2C03
        "--------", -- 0x2C04
        "--------", -- 0x2C05
        "--------", -- 0x2C06
        "--------", -- 0x2C07
        "--------", -- 0x2C08
        "--------", -- 0x2C09
        "--------", -- 0x2C0A
        "--------", -- 0x2C0B
        "--------", -- 0x2C0C
        "--------", -- 0x2C0D
        "--------", -- 0x2C0E
        "--------", -- 0x2C0F
        "--------", -- 0x2C10
        "--------", -- 0x2C11
        "--------", -- 0x2C12
        "--------", -- 0x2C13
        "--------", -- 0x2C14
        "--------", -- 0x2C15
        "--------", -- 0x2C16
        "--------", -- 0x2C17
        "--------", -- 0x2C18
        "--------", -- 0x2C19
        "--------", -- 0x2C1A
        "--------", -- 0x2C1B
        "--------", -- 0x2C1C
        "--------", -- 0x2C1D
        "--------", -- 0x2C1E
        "--------", -- 0x2C1F
        "--------", -- 0x2C20
        "--------", -- 0x2C21
        "--------", -- 0x2C22
        "--------", -- 0x2C23
        "--------", -- 0x2C24
        "--------", -- 0x2C25
        "--------", -- 0x2C26
        "--------", -- 0x2C27
        "--------", -- 0x2C28
        "--------", -- 0x2C29
        "--------", -- 0x2C2A
        "--------", -- 0x2C2B
        "--------", -- 0x2C2C
        "--------", -- 0x2C2D
        "--------", -- 0x2C2E
        "--------", -- 0x2C2F
        "--------", -- 0x2C30
        "--------", -- 0x2C31
        "--------", -- 0x2C32
        "--------", -- 0x2C33
        "--------", -- 0x2C34
        "--------", -- 0x2C35
        "--------", -- 0x2C36
        "--------", -- 0x2C37
        "--------", -- 0x2C38
        "--------", -- 0x2C39
        "--------", -- 0x2C3A
        "--------", -- 0x2C3B
        "--------", -- 0x2C3C
        "--------", -- 0x2C3D
        "--------", -- 0x2C3E
        "--------", -- 0x2C3F
        "--------", -- 0x2C40
        "--------", -- 0x2C41
        "--------", -- 0x2C42
        "--------", -- 0x2C43
        "--------", -- 0x2C44
        "--------", -- 0x2C45
        "--------", -- 0x2C46
        "--------", -- 0x2C47
        "--------", -- 0x2C48
        "--------", -- 0x2C49
        "--------", -- 0x2C4A
        "--------", -- 0x2C4B
        "--------", -- 0x2C4C
        "--------", -- 0x2C4D
        "--------", -- 0x2C4E
        "--------", -- 0x2C4F
        "--------", -- 0x2C50
        "--------", -- 0x2C51
        "--------", -- 0x2C52
        "--------", -- 0x2C53
        "--------", -- 0x2C54
        "--------", -- 0x2C55
        "--------", -- 0x2C56
        "--------", -- 0x2C57
        "--------", -- 0x2C58
        "--------", -- 0x2C59
        "--------", -- 0x2C5A
        "--------", -- 0x2C5B
        "--------", -- 0x2C5C
        "--------", -- 0x2C5D
        "--------", -- 0x2C5E
        "--------", -- 0x2C5F
        "--------", -- 0x2C60
        "--------", -- 0x2C61
        "--------", -- 0x2C62
        "--------", -- 0x2C63
        "--------", -- 0x2C64
        "--------", -- 0x2C65
        "--------", -- 0x2C66
        "--------", -- 0x2C67
        "--------", -- 0x2C68
        "--------", -- 0x2C69
        "--------", -- 0x2C6A
        "--------", -- 0x2C6B
        "--------", -- 0x2C6C
        "--------", -- 0x2C6D
        "--------", -- 0x2C6E
        "--------", -- 0x2C6F
        "--------", -- 0x2C70
        "--------", -- 0x2C71
        "--------", -- 0x2C72
        "--------", -- 0x2C73
        "--------", -- 0x2C74
        "--------", -- 0x2C75
        "--------", -- 0x2C76
        "--------", -- 0x2C77
        "--------", -- 0x2C78
        "--------", -- 0x2C79
        "--------", -- 0x2C7A
        "--------", -- 0x2C7B
        "--------", -- 0x2C7C
        "--------", -- 0x2C7D
        "--------", -- 0x2C7E
        "--------", -- 0x2C7F
        "--------", -- 0x2C80
        "--------", -- 0x2C81
        "--------", -- 0x2C82
        "--------", -- 0x2C83
        "--------", -- 0x2C84
        "--------", -- 0x2C85
        "--------", -- 0x2C86
        "--------", -- 0x2C87
        "--------", -- 0x2C88
        "--------", -- 0x2C89
        "--------", -- 0x2C8A
        "--------", -- 0x2C8B
        "--------", -- 0x2C8C
        "--------", -- 0x2C8D
        "--------", -- 0x2C8E
        "--------", -- 0x2C8F
        "--------", -- 0x2C90
        "--------", -- 0x2C91
        "--------", -- 0x2C92
        "--------", -- 0x2C93
        "--------", -- 0x2C94
        "--------", -- 0x2C95
        "--------", -- 0x2C96
        "--------", -- 0x2C97
        "--------", -- 0x2C98
        "--------", -- 0x2C99
        "--------", -- 0x2C9A
        "--------", -- 0x2C9B
        "--------", -- 0x2C9C
        "--------", -- 0x2C9D
        "--------", -- 0x2C9E
        "--------", -- 0x2C9F
        "--------", -- 0x2CA0
        "--------", -- 0x2CA1
        "--------", -- 0x2CA2
        "--------", -- 0x2CA3
        "--------", -- 0x2CA4
        "--------", -- 0x2CA5
        "--------", -- 0x2CA6
        "--------", -- 0x2CA7
        "--------", -- 0x2CA8
        "--------", -- 0x2CA9
        "--------", -- 0x2CAA
        "--------", -- 0x2CAB
        "--------", -- 0x2CAC
        "--------", -- 0x2CAD
        "--------", -- 0x2CAE
        "--------", -- 0x2CAF
        "--------", -- 0x2CB0
        "--------", -- 0x2CB1
        "--------", -- 0x2CB2
        "--------", -- 0x2CB3
        "--------", -- 0x2CB4
        "--------", -- 0x2CB5
        "--------", -- 0x2CB6
        "--------", -- 0x2CB7
        "--------", -- 0x2CB8
        "--------", -- 0x2CB9
        "--------", -- 0x2CBA
        "--------", -- 0x2CBB
        "--------", -- 0x2CBC
        "--------", -- 0x2CBD
        "--------", -- 0x2CBE
        "--------", -- 0x2CBF
        "--------", -- 0x2CC0
        "--------", -- 0x2CC1
        "--------", -- 0x2CC2
        "--------", -- 0x2CC3
        "--------", -- 0x2CC4
        "--------", -- 0x2CC5
        "--------", -- 0x2CC6
        "--------", -- 0x2CC7
        "--------", -- 0x2CC8
        "--------", -- 0x2CC9
        "--------", -- 0x2CCA
        "--------", -- 0x2CCB
        "--------", -- 0x2CCC
        "--------", -- 0x2CCD
        "--------", -- 0x2CCE
        "--------", -- 0x2CCF
        "--------", -- 0x2CD0
        "--------", -- 0x2CD1
        "--------", -- 0x2CD2
        "--------", -- 0x2CD3
        "--------", -- 0x2CD4
        "--------", -- 0x2CD5
        "--------", -- 0x2CD6
        "--------", -- 0x2CD7
        "--------", -- 0x2CD8
        "--------", -- 0x2CD9
        "--------", -- 0x2CDA
        "--------", -- 0x2CDB
        "--------", -- 0x2CDC
        "--------", -- 0x2CDD
        "--------", -- 0x2CDE
        "--------", -- 0x2CDF
        "--------", -- 0x2CE0
        "--------", -- 0x2CE1
        "--------", -- 0x2CE2
        "--------", -- 0x2CE3
        "--------", -- 0x2CE4
        "--------", -- 0x2CE5
        "--------", -- 0x2CE6
        "--------", -- 0x2CE7
        "--------", -- 0x2CE8
        "--------", -- 0x2CE9
        "--------", -- 0x2CEA
        "--------", -- 0x2CEB
        "--------", -- 0x2CEC
        "--------", -- 0x2CED
        "--------", -- 0x2CEE
        "--------", -- 0x2CEF
        "--------", -- 0x2CF0
        "--------", -- 0x2CF1
        "--------", -- 0x2CF2
        "--------", -- 0x2CF3
        "--------", -- 0x2CF4
        "--------", -- 0x2CF5
        "--------", -- 0x2CF6
        "--------", -- 0x2CF7
        "--------", -- 0x2CF8
        "--------", -- 0x2CF9
        "--------", -- 0x2CFA
        "--------", -- 0x2CFB
        "--------", -- 0x2CFC
        "--------", -- 0x2CFD
        "--------", -- 0x2CFE
        "--------", -- 0x2CFF
        "--------", -- 0x2D00
        "--------", -- 0x2D01
        "--------", -- 0x2D02
        "--------", -- 0x2D03
        "--------", -- 0x2D04
        "--------", -- 0x2D05
        "--------", -- 0x2D06
        "--------", -- 0x2D07
        "--------", -- 0x2D08
        "--------", -- 0x2D09
        "--------", -- 0x2D0A
        "--------", -- 0x2D0B
        "--------", -- 0x2D0C
        "--------", -- 0x2D0D
        "--------", -- 0x2D0E
        "--------", -- 0x2D0F
        "--------", -- 0x2D10
        "--------", -- 0x2D11
        "--------", -- 0x2D12
        "--------", -- 0x2D13
        "--------", -- 0x2D14
        "--------", -- 0x2D15
        "--------", -- 0x2D16
        "--------", -- 0x2D17
        "--------", -- 0x2D18
        "--------", -- 0x2D19
        "--------", -- 0x2D1A
        "--------", -- 0x2D1B
        "--------", -- 0x2D1C
        "--------", -- 0x2D1D
        "--------", -- 0x2D1E
        "--------", -- 0x2D1F
        "--------", -- 0x2D20
        "--------", -- 0x2D21
        "--------", -- 0x2D22
        "--------", -- 0x2D23
        "--------", -- 0x2D24
        "--------", -- 0x2D25
        "--------", -- 0x2D26
        "--------", -- 0x2D27
        "--------", -- 0x2D28
        "--------", -- 0x2D29
        "--------", -- 0x2D2A
        "--------", -- 0x2D2B
        "--------", -- 0x2D2C
        "--------", -- 0x2D2D
        "--------", -- 0x2D2E
        "--------", -- 0x2D2F
        "--------", -- 0x2D30
        "--------", -- 0x2D31
        "--------", -- 0x2D32
        "--------", -- 0x2D33
        "--------", -- 0x2D34
        "--------", -- 0x2D35
        "--------", -- 0x2D36
        "--------", -- 0x2D37
        "--------", -- 0x2D38
        "--------", -- 0x2D39
        "--------", -- 0x2D3A
        "--------", -- 0x2D3B
        "--------", -- 0x2D3C
        "--------", -- 0x2D3D
        "--------", -- 0x2D3E
        "--------", -- 0x2D3F
        "--------", -- 0x2D40
        "--------", -- 0x2D41
        "--------", -- 0x2D42
        "--------", -- 0x2D43
        "--------", -- 0x2D44
        "--------", -- 0x2D45
        "--------", -- 0x2D46
        "--------", -- 0x2D47
        "--------", -- 0x2D48
        "--------", -- 0x2D49
        "--------", -- 0x2D4A
        "--------", -- 0x2D4B
        "--------", -- 0x2D4C
        "--------", -- 0x2D4D
        "--------", -- 0x2D4E
        "--------", -- 0x2D4F
        "--------", -- 0x2D50
        "--------", -- 0x2D51
        "--------", -- 0x2D52
        "--------", -- 0x2D53
        "--------", -- 0x2D54
        "--------", -- 0x2D55
        "--------", -- 0x2D56
        "--------", -- 0x2D57
        "--------", -- 0x2D58
        "--------", -- 0x2D59
        "--------", -- 0x2D5A
        "--------", -- 0x2D5B
        "--------", -- 0x2D5C
        "--------", -- 0x2D5D
        "--------", -- 0x2D5E
        "--------", -- 0x2D5F
        "--------", -- 0x2D60
        "--------", -- 0x2D61
        "--------", -- 0x2D62
        "--------", -- 0x2D63
        "--------", -- 0x2D64
        "--------", -- 0x2D65
        "--------", -- 0x2D66
        "--------", -- 0x2D67
        "--------", -- 0x2D68
        "--------", -- 0x2D69
        "--------", -- 0x2D6A
        "--------", -- 0x2D6B
        "--------", -- 0x2D6C
        "--------", -- 0x2D6D
        "--------", -- 0x2D6E
        "--------", -- 0x2D6F
        "--------", -- 0x2D70
        "--------", -- 0x2D71
        "--------", -- 0x2D72
        "--------", -- 0x2D73
        "--------", -- 0x2D74
        "--------", -- 0x2D75
        "--------", -- 0x2D76
        "--------", -- 0x2D77
        "--------", -- 0x2D78
        "--------", -- 0x2D79
        "--------", -- 0x2D7A
        "--------", -- 0x2D7B
        "--------", -- 0x2D7C
        "--------", -- 0x2D7D
        "--------", -- 0x2D7E
        "--------", -- 0x2D7F
        "--------", -- 0x2D80
        "--------", -- 0x2D81
        "--------", -- 0x2D82
        "--------", -- 0x2D83
        "--------", -- 0x2D84
        "--------", -- 0x2D85
        "--------", -- 0x2D86
        "--------", -- 0x2D87
        "--------", -- 0x2D88
        "--------", -- 0x2D89
        "--------", -- 0x2D8A
        "--------", -- 0x2D8B
        "--------", -- 0x2D8C
        "--------", -- 0x2D8D
        "--------", -- 0x2D8E
        "--------", -- 0x2D8F
        "--------", -- 0x2D90
        "--------", -- 0x2D91
        "--------", -- 0x2D92
        "--------", -- 0x2D93
        "--------", -- 0x2D94
        "--------", -- 0x2D95
        "--------", -- 0x2D96
        "--------", -- 0x2D97
        "--------", -- 0x2D98
        "--------", -- 0x2D99
        "--------", -- 0x2D9A
        "--------", -- 0x2D9B
        "--------", -- 0x2D9C
        "--------", -- 0x2D9D
        "--------", -- 0x2D9E
        "--------", -- 0x2D9F
        "--------", -- 0x2DA0
        "--------", -- 0x2DA1
        "--------", -- 0x2DA2
        "--------", -- 0x2DA3
        "--------", -- 0x2DA4
        "--------", -- 0x2DA5
        "--------", -- 0x2DA6
        "--------", -- 0x2DA7
        "--------", -- 0x2DA8
        "--------", -- 0x2DA9
        "--------", -- 0x2DAA
        "--------", -- 0x2DAB
        "--------", -- 0x2DAC
        "--------", -- 0x2DAD
        "--------", -- 0x2DAE
        "--------", -- 0x2DAF
        "--------", -- 0x2DB0
        "--------", -- 0x2DB1
        "--------", -- 0x2DB2
        "--------", -- 0x2DB3
        "--------", -- 0x2DB4
        "--------", -- 0x2DB5
        "--------", -- 0x2DB6
        "--------", -- 0x2DB7
        "--------", -- 0x2DB8
        "--------", -- 0x2DB9
        "--------", -- 0x2DBA
        "--------", -- 0x2DBB
        "--------", -- 0x2DBC
        "--------", -- 0x2DBD
        "--------", -- 0x2DBE
        "--------", -- 0x2DBF
        "--------", -- 0x2DC0
        "--------", -- 0x2DC1
        "--------", -- 0x2DC2
        "--------", -- 0x2DC3
        "--------", -- 0x2DC4
        "--------", -- 0x2DC5
        "--------", -- 0x2DC6
        "--------", -- 0x2DC7
        "--------", -- 0x2DC8
        "--------", -- 0x2DC9
        "--------", -- 0x2DCA
        "--------", -- 0x2DCB
        "--------", -- 0x2DCC
        "--------", -- 0x2DCD
        "--------", -- 0x2DCE
        "--------", -- 0x2DCF
        "--------", -- 0x2DD0
        "--------", -- 0x2DD1
        "--------", -- 0x2DD2
        "--------", -- 0x2DD3
        "--------", -- 0x2DD4
        "--------", -- 0x2DD5
        "--------", -- 0x2DD6
        "--------", -- 0x2DD7
        "--------", -- 0x2DD8
        "--------", -- 0x2DD9
        "--------", -- 0x2DDA
        "--------", -- 0x2DDB
        "--------", -- 0x2DDC
        "--------", -- 0x2DDD
        "--------", -- 0x2DDE
        "--------", -- 0x2DDF
        "--------", -- 0x2DE0
        "--------", -- 0x2DE1
        "--------", -- 0x2DE2
        "--------", -- 0x2DE3
        "--------", -- 0x2DE4
        "--------", -- 0x2DE5
        "--------", -- 0x2DE6
        "--------", -- 0x2DE7
        "--------", -- 0x2DE8
        "--------", -- 0x2DE9
        "--------", -- 0x2DEA
        "--------", -- 0x2DEB
        "--------", -- 0x2DEC
        "--------", -- 0x2DED
        "--------", -- 0x2DEE
        "--------", -- 0x2DEF
        "--------", -- 0x2DF0
        "--------", -- 0x2DF1
        "--------", -- 0x2DF2
        "--------", -- 0x2DF3
        "--------", -- 0x2DF4
        "--------", -- 0x2DF5
        "--------", -- 0x2DF6
        "--------", -- 0x2DF7
        "--------", -- 0x2DF8
        "--------", -- 0x2DF9
        "--------", -- 0x2DFA
        "--------", -- 0x2DFB
        "--------", -- 0x2DFC
        "--------", -- 0x2DFD
        "--------", -- 0x2DFE
        "--------", -- 0x2DFF
        "--------", -- 0x2E00
        "--------", -- 0x2E01
        "--------", -- 0x2E02
        "--------", -- 0x2E03
        "--------", -- 0x2E04
        "--------", -- 0x2E05
        "--------", -- 0x2E06
        "--------", -- 0x2E07
        "--------", -- 0x2E08
        "--------", -- 0x2E09
        "--------", -- 0x2E0A
        "--------", -- 0x2E0B
        "--------", -- 0x2E0C
        "--------", -- 0x2E0D
        "--------", -- 0x2E0E
        "--------", -- 0x2E0F
        "--------", -- 0x2E10
        "--------", -- 0x2E11
        "--------", -- 0x2E12
        "--------", -- 0x2E13
        "--------", -- 0x2E14
        "--------", -- 0x2E15
        "--------", -- 0x2E16
        "--------", -- 0x2E17
        "--------", -- 0x2E18
        "--------", -- 0x2E19
        "--------", -- 0x2E1A
        "--------", -- 0x2E1B
        "--------", -- 0x2E1C
        "--------", -- 0x2E1D
        "--------", -- 0x2E1E
        "--------", -- 0x2E1F
        "--------", -- 0x2E20
        "--------", -- 0x2E21
        "--------", -- 0x2E22
        "--------", -- 0x2E23
        "--------", -- 0x2E24
        "--------", -- 0x2E25
        "--------", -- 0x2E26
        "--------", -- 0x2E27
        "--------", -- 0x2E28
        "--------", -- 0x2E29
        "--------", -- 0x2E2A
        "--------", -- 0x2E2B
        "--------", -- 0x2E2C
        "--------", -- 0x2E2D
        "--------", -- 0x2E2E
        "--------", -- 0x2E2F
        "--------", -- 0x2E30
        "--------", -- 0x2E31
        "--------", -- 0x2E32
        "--------", -- 0x2E33
        "--------", -- 0x2E34
        "--------", -- 0x2E35
        "--------", -- 0x2E36
        "--------", -- 0x2E37
        "--------", -- 0x2E38
        "--------", -- 0x2E39
        "--------", -- 0x2E3A
        "--------", -- 0x2E3B
        "--------", -- 0x2E3C
        "--------", -- 0x2E3D
        "--------", -- 0x2E3E
        "--------", -- 0x2E3F
        "--------", -- 0x2E40
        "--------", -- 0x2E41
        "--------", -- 0x2E42
        "--------", -- 0x2E43
        "--------", -- 0x2E44
        "--------", -- 0x2E45
        "--------", -- 0x2E46
        "--------", -- 0x2E47
        "--------", -- 0x2E48
        "--------", -- 0x2E49
        "--------", -- 0x2E4A
        "--------", -- 0x2E4B
        "--------", -- 0x2E4C
        "--------", -- 0x2E4D
        "--------", -- 0x2E4E
        "--------", -- 0x2E4F
        "--------", -- 0x2E50
        "--------", -- 0x2E51
        "--------", -- 0x2E52
        "--------", -- 0x2E53
        "--------", -- 0x2E54
        "--------", -- 0x2E55
        "--------", -- 0x2E56
        "--------", -- 0x2E57
        "--------", -- 0x2E58
        "--------", -- 0x2E59
        "--------", -- 0x2E5A
        "--------", -- 0x2E5B
        "--------", -- 0x2E5C
        "--------", -- 0x2E5D
        "--------", -- 0x2E5E
        "--------", -- 0x2E5F
        "--------", -- 0x2E60
        "--------", -- 0x2E61
        "--------", -- 0x2E62
        "--------", -- 0x2E63
        "--------", -- 0x2E64
        "--------", -- 0x2E65
        "--------", -- 0x2E66
        "--------", -- 0x2E67
        "--------", -- 0x2E68
        "--------", -- 0x2E69
        "--------", -- 0x2E6A
        "--------", -- 0x2E6B
        "--------", -- 0x2E6C
        "--------", -- 0x2E6D
        "--------", -- 0x2E6E
        "--------", -- 0x2E6F
        "--------", -- 0x2E70
        "--------", -- 0x2E71
        "--------", -- 0x2E72
        "--------", -- 0x2E73
        "--------", -- 0x2E74
        "--------", -- 0x2E75
        "--------", -- 0x2E76
        "--------", -- 0x2E77
        "--------", -- 0x2E78
        "--------", -- 0x2E79
        "--------", -- 0x2E7A
        "--------", -- 0x2E7B
        "--------", -- 0x2E7C
        "--------", -- 0x2E7D
        "--------", -- 0x2E7E
        "--------", -- 0x2E7F
        "--------", -- 0x2E80
        "--------", -- 0x2E81
        "--------", -- 0x2E82
        "--------", -- 0x2E83
        "--------", -- 0x2E84
        "--------", -- 0x2E85
        "--------", -- 0x2E86
        "--------", -- 0x2E87
        "--------", -- 0x2E88
        "--------", -- 0x2E89
        "--------", -- 0x2E8A
        "--------", -- 0x2E8B
        "--------", -- 0x2E8C
        "--------", -- 0x2E8D
        "--------", -- 0x2E8E
        "--------", -- 0x2E8F
        "--------", -- 0x2E90
        "--------", -- 0x2E91
        "--------", -- 0x2E92
        "--------", -- 0x2E93
        "--------", -- 0x2E94
        "--------", -- 0x2E95
        "--------", -- 0x2E96
        "--------", -- 0x2E97
        "--------", -- 0x2E98
        "--------", -- 0x2E99
        "--------", -- 0x2E9A
        "--------", -- 0x2E9B
        "--------", -- 0x2E9C
        "--------", -- 0x2E9D
        "--------", -- 0x2E9E
        "--------", -- 0x2E9F
        "--------", -- 0x2EA0
        "--------", -- 0x2EA1
        "--------", -- 0x2EA2
        "--------", -- 0x2EA3
        "--------", -- 0x2EA4
        "--------", -- 0x2EA5
        "--------", -- 0x2EA6
        "--------", -- 0x2EA7
        "--------", -- 0x2EA8
        "--------", -- 0x2EA9
        "--------", -- 0x2EAA
        "--------", -- 0x2EAB
        "--------", -- 0x2EAC
        "--------", -- 0x2EAD
        "--------", -- 0x2EAE
        "--------", -- 0x2EAF
        "--------", -- 0x2EB0
        "--------", -- 0x2EB1
        "--------", -- 0x2EB2
        "--------", -- 0x2EB3
        "--------", -- 0x2EB4
        "--------", -- 0x2EB5
        "--------", -- 0x2EB6
        "--------", -- 0x2EB7
        "--------", -- 0x2EB8
        "--------", -- 0x2EB9
        "--------", -- 0x2EBA
        "--------", -- 0x2EBB
        "--------", -- 0x2EBC
        "--------", -- 0x2EBD
        "--------", -- 0x2EBE
        "--------", -- 0x2EBF
        "--------", -- 0x2EC0
        "--------", -- 0x2EC1
        "--------", -- 0x2EC2
        "--------", -- 0x2EC3
        "--------", -- 0x2EC4
        "--------", -- 0x2EC5
        "--------", -- 0x2EC6
        "--------", -- 0x2EC7
        "--------", -- 0x2EC8
        "--------", -- 0x2EC9
        "--------", -- 0x2ECA
        "--------", -- 0x2ECB
        "--------", -- 0x2ECC
        "--------", -- 0x2ECD
        "--------", -- 0x2ECE
        "--------", -- 0x2ECF
        "--------", -- 0x2ED0
        "--------", -- 0x2ED1
        "--------", -- 0x2ED2
        "--------", -- 0x2ED3
        "--------", -- 0x2ED4
        "--------", -- 0x2ED5
        "--------", -- 0x2ED6
        "--------", -- 0x2ED7
        "--------", -- 0x2ED8
        "--------", -- 0x2ED9
        "--------", -- 0x2EDA
        "--------", -- 0x2EDB
        "--------", -- 0x2EDC
        "--------", -- 0x2EDD
        "--------", -- 0x2EDE
        "--------", -- 0x2EDF
        "--------", -- 0x2EE0
        "--------", -- 0x2EE1
        "--------", -- 0x2EE2
        "--------", -- 0x2EE3
        "--------", -- 0x2EE4
        "--------", -- 0x2EE5
        "--------", -- 0x2EE6
        "--------", -- 0x2EE7
        "--------", -- 0x2EE8
        "--------", -- 0x2EE9
        "--------", -- 0x2EEA
        "--------", -- 0x2EEB
        "--------", -- 0x2EEC
        "--------", -- 0x2EED
        "--------", -- 0x2EEE
        "--------", -- 0x2EEF
        "--------", -- 0x2EF0
        "--------", -- 0x2EF1
        "--------", -- 0x2EF2
        "--------", -- 0x2EF3
        "--------", -- 0x2EF4
        "--------", -- 0x2EF5
        "--------", -- 0x2EF6
        "--------", -- 0x2EF7
        "--------", -- 0x2EF8
        "--------", -- 0x2EF9
        "--------", -- 0x2EFA
        "--------", -- 0x2EFB
        "--------", -- 0x2EFC
        "--------", -- 0x2EFD
        "--------", -- 0x2EFE
        "--------", -- 0x2EFF
        "--------", -- 0x2F00
        "--------", -- 0x2F01
        "--------", -- 0x2F02
        "--------", -- 0x2F03
        "--------", -- 0x2F04
        "--------", -- 0x2F05
        "--------", -- 0x2F06
        "--------", -- 0x2F07
        "--------", -- 0x2F08
        "--------", -- 0x2F09
        "--------", -- 0x2F0A
        "--------", -- 0x2F0B
        "--------", -- 0x2F0C
        "--------", -- 0x2F0D
        "--------", -- 0x2F0E
        "--------", -- 0x2F0F
        "--------", -- 0x2F10
        "--------", -- 0x2F11
        "--------", -- 0x2F12
        "--------", -- 0x2F13
        "--------", -- 0x2F14
        "--------", -- 0x2F15
        "--------", -- 0x2F16
        "--------", -- 0x2F17
        "--------", -- 0x2F18
        "--------", -- 0x2F19
        "--------", -- 0x2F1A
        "--------", -- 0x2F1B
        "--------", -- 0x2F1C
        "--------", -- 0x2F1D
        "--------", -- 0x2F1E
        "--------", -- 0x2F1F
        "--------", -- 0x2F20
        "--------", -- 0x2F21
        "--------", -- 0x2F22
        "--------", -- 0x2F23
        "--------", -- 0x2F24
        "--------", -- 0x2F25
        "--------", -- 0x2F26
        "--------", -- 0x2F27
        "--------", -- 0x2F28
        "--------", -- 0x2F29
        "--------", -- 0x2F2A
        "--------", -- 0x2F2B
        "--------", -- 0x2F2C
        "--------", -- 0x2F2D
        "--------", -- 0x2F2E
        "--------", -- 0x2F2F
        "--------", -- 0x2F30
        "--------", -- 0x2F31
        "--------", -- 0x2F32
        "--------", -- 0x2F33
        "--------", -- 0x2F34
        "--------", -- 0x2F35
        "--------", -- 0x2F36
        "--------", -- 0x2F37
        "--------", -- 0x2F38
        "--------", -- 0x2F39
        "--------", -- 0x2F3A
        "--------", -- 0x2F3B
        "--------", -- 0x2F3C
        "--------", -- 0x2F3D
        "--------", -- 0x2F3E
        "--------", -- 0x2F3F
        "--------", -- 0x2F40
        "--------", -- 0x2F41
        "--------", -- 0x2F42
        "--------", -- 0x2F43
        "--------", -- 0x2F44
        "--------", -- 0x2F45
        "--------", -- 0x2F46
        "--------", -- 0x2F47
        "--------", -- 0x2F48
        "--------", -- 0x2F49
        "--------", -- 0x2F4A
        "--------", -- 0x2F4B
        "--------", -- 0x2F4C
        "--------", -- 0x2F4D
        "--------", -- 0x2F4E
        "--------", -- 0x2F4F
        "--------", -- 0x2F50
        "--------", -- 0x2F51
        "--------", -- 0x2F52
        "--------", -- 0x2F53
        "--------", -- 0x2F54
        "--------", -- 0x2F55
        "--------", -- 0x2F56
        "--------", -- 0x2F57
        "--------", -- 0x2F58
        "--------", -- 0x2F59
        "--------", -- 0x2F5A
        "--------", -- 0x2F5B
        "--------", -- 0x2F5C
        "--------", -- 0x2F5D
        "--------", -- 0x2F5E
        "--------", -- 0x2F5F
        "--------", -- 0x2F60
        "--------", -- 0x2F61
        "--------", -- 0x2F62
        "--------", -- 0x2F63
        "--------", -- 0x2F64
        "--------", -- 0x2F65
        "--------", -- 0x2F66
        "--------", -- 0x2F67
        "--------", -- 0x2F68
        "--------", -- 0x2F69
        "--------", -- 0x2F6A
        "--------", -- 0x2F6B
        "--------", -- 0x2F6C
        "--------", -- 0x2F6D
        "--------", -- 0x2F6E
        "--------", -- 0x2F6F
        "--------", -- 0x2F70
        "--------", -- 0x2F71
        "--------", -- 0x2F72
        "--------", -- 0x2F73
        "--------", -- 0x2F74
        "--------", -- 0x2F75
        "--------", -- 0x2F76
        "--------", -- 0x2F77
        "--------", -- 0x2F78
        "--------", -- 0x2F79
        "--------", -- 0x2F7A
        "--------", -- 0x2F7B
        "--------", -- 0x2F7C
        "--------", -- 0x2F7D
        "--------", -- 0x2F7E
        "--------", -- 0x2F7F
        "--------", -- 0x2F80
        "--------", -- 0x2F81
        "--------", -- 0x2F82
        "--------", -- 0x2F83
        "--------", -- 0x2F84
        "--------", -- 0x2F85
        "--------", -- 0x2F86
        "--------", -- 0x2F87
        "--------", -- 0x2F88
        "--------", -- 0x2F89
        "--------", -- 0x2F8A
        "--------", -- 0x2F8B
        "--------", -- 0x2F8C
        "--------", -- 0x2F8D
        "--------", -- 0x2F8E
        "--------", -- 0x2F8F
        "--------", -- 0x2F90
        "--------", -- 0x2F91
        "--------", -- 0x2F92
        "--------", -- 0x2F93
        "--------", -- 0x2F94
        "--------", -- 0x2F95
        "--------", -- 0x2F96
        "--------", -- 0x2F97
        "--------", -- 0x2F98
        "--------", -- 0x2F99
        "--------", -- 0x2F9A
        "--------", -- 0x2F9B
        "--------", -- 0x2F9C
        "--------", -- 0x2F9D
        "--------", -- 0x2F9E
        "--------", -- 0x2F9F
        "--------", -- 0x2FA0
        "--------", -- 0x2FA1
        "--------", -- 0x2FA2
        "--------", -- 0x2FA3
        "--------", -- 0x2FA4
        "--------", -- 0x2FA5
        "--------", -- 0x2FA6
        "--------", -- 0x2FA7
        "--------", -- 0x2FA8
        "--------", -- 0x2FA9
        "--------", -- 0x2FAA
        "--------", -- 0x2FAB
        "--------", -- 0x2FAC
        "--------", -- 0x2FAD
        "--------", -- 0x2FAE
        "--------", -- 0x2FAF
        "--------", -- 0x2FB0
        "--------", -- 0x2FB1
        "--------", -- 0x2FB2
        "--------", -- 0x2FB3
        "--------", -- 0x2FB4
        "--------", -- 0x2FB5
        "--------", -- 0x2FB6
        "--------", -- 0x2FB7
        "--------", -- 0x2FB8
        "--------", -- 0x2FB9
        "--------", -- 0x2FBA
        "--------", -- 0x2FBB
        "--------", -- 0x2FBC
        "--------", -- 0x2FBD
        "--------", -- 0x2FBE
        "--------", -- 0x2FBF
        "--------", -- 0x2FC0
        "--------", -- 0x2FC1
        "--------", -- 0x2FC2
        "--------", -- 0x2FC3
        "--------", -- 0x2FC4
        "--------", -- 0x2FC5
        "--------", -- 0x2FC6
        "--------", -- 0x2FC7
        "--------", -- 0x2FC8
        "--------", -- 0x2FC9
        "--------", -- 0x2FCA
        "--------", -- 0x2FCB
        "--------", -- 0x2FCC
        "--------", -- 0x2FCD
        "--------", -- 0x2FCE
        "--------", -- 0x2FCF
        "--------", -- 0x2FD0
        "--------", -- 0x2FD1
        "--------", -- 0x2FD2
        "--------", -- 0x2FD3
        "--------", -- 0x2FD4
        "--------", -- 0x2FD5
        "--------", -- 0x2FD6
        "--------", -- 0x2FD7
        "--------", -- 0x2FD8
        "--------", -- 0x2FD9
        "--------", -- 0x2FDA
        "--------", -- 0x2FDB
        "--------", -- 0x2FDC
        "--------", -- 0x2FDD
        "--------", -- 0x2FDE
        "--------", -- 0x2FDF
        "--------", -- 0x2FE0
        "--------", -- 0x2FE1
        "--------", -- 0x2FE2
        "--------", -- 0x2FE3
        "--------", -- 0x2FE4
        "--------", -- 0x2FE5
        "--------", -- 0x2FE6
        "--------", -- 0x2FE7
        "--------", -- 0x2FE8
        "--------", -- 0x2FE9
        "--------", -- 0x2FEA
        "--------", -- 0x2FEB
        "--------", -- 0x2FEC
        "--------", -- 0x2FED
        "--------", -- 0x2FEE
        "--------", -- 0x2FEF
        "--------", -- 0x2FF0
        "--------", -- 0x2FF1
        "--------", -- 0x2FF2
        "--------", -- 0x2FF3
        "--------", -- 0x2FF4
        "--------", -- 0x2FF5
        "--------", -- 0x2FF6
        "--------", -- 0x2FF7
        "--------", -- 0x2FF8
        "--------", -- 0x2FF9
        "--------", -- 0x2FFA
        "--------", -- 0x2FFB
        "--------", -- 0x2FFC
        "--------", -- 0x2FFD
        "--------", -- 0x2FFE
        "--------", -- 0x2FFF
        "--------", -- 0x3000
        "--------", -- 0x3001
        "--------", -- 0x3002
        "--------", -- 0x3003
        "--------", -- 0x3004
        "--------", -- 0x3005
        "--------", -- 0x3006
        "--------", -- 0x3007
        "--------", -- 0x3008
        "--------", -- 0x3009
        "--------", -- 0x300A
        "--------", -- 0x300B
        "--------", -- 0x300C
        "--------", -- 0x300D
        "--------", -- 0x300E
        "--------", -- 0x300F
        "--------", -- 0x3010
        "--------", -- 0x3011
        "--------", -- 0x3012
        "--------", -- 0x3013
        "--------", -- 0x3014
        "--------", -- 0x3015
        "--------", -- 0x3016
        "--------", -- 0x3017
        "--------", -- 0x3018
        "--------", -- 0x3019
        "--------", -- 0x301A
        "--------", -- 0x301B
        "--------", -- 0x301C
        "--------", -- 0x301D
        "--------", -- 0x301E
        "--------", -- 0x301F
        "--------", -- 0x3020
        "--------", -- 0x3021
        "--------", -- 0x3022
        "--------", -- 0x3023
        "--------", -- 0x3024
        "--------", -- 0x3025
        "--------", -- 0x3026
        "--------", -- 0x3027
        "--------", -- 0x3028
        "--------", -- 0x3029
        "--------", -- 0x302A
        "--------", -- 0x302B
        "--------", -- 0x302C
        "--------", -- 0x302D
        "--------", -- 0x302E
        "--------", -- 0x302F
        "--------", -- 0x3030
        "--------", -- 0x3031
        "--------", -- 0x3032
        "--------", -- 0x3033
        "--------", -- 0x3034
        "--------", -- 0x3035
        "--------", -- 0x3036
        "--------", -- 0x3037
        "--------", -- 0x3038
        "--------", -- 0x3039
        "--------", -- 0x303A
        "--------", -- 0x303B
        "--------", -- 0x303C
        "--------", -- 0x303D
        "--------", -- 0x303E
        "--------", -- 0x303F
        "--------", -- 0x3040
        "--------", -- 0x3041
        "--------", -- 0x3042
        "--------", -- 0x3043
        "--------", -- 0x3044
        "--------", -- 0x3045
        "--------", -- 0x3046
        "--------", -- 0x3047
        "--------", -- 0x3048
        "--------", -- 0x3049
        "--------", -- 0x304A
        "--------", -- 0x304B
        "--------", -- 0x304C
        "--------", -- 0x304D
        "--------", -- 0x304E
        "--------", -- 0x304F
        "--------", -- 0x3050
        "--------", -- 0x3051
        "--------", -- 0x3052
        "--------", -- 0x3053
        "--------", -- 0x3054
        "--------", -- 0x3055
        "--------", -- 0x3056
        "--------", -- 0x3057
        "--------", -- 0x3058
        "--------", -- 0x3059
        "--------", -- 0x305A
        "--------", -- 0x305B
        "--------", -- 0x305C
        "--------", -- 0x305D
        "--------", -- 0x305E
        "--------", -- 0x305F
        "--------", -- 0x3060
        "--------", -- 0x3061
        "--------", -- 0x3062
        "--------", -- 0x3063
        "--------", -- 0x3064
        "--------", -- 0x3065
        "--------", -- 0x3066
        "--------", -- 0x3067
        "--------", -- 0x3068
        "--------", -- 0x3069
        "--------", -- 0x306A
        "--------", -- 0x306B
        "--------", -- 0x306C
        "--------", -- 0x306D
        "--------", -- 0x306E
        "--------", -- 0x306F
        "--------", -- 0x3070
        "--------", -- 0x3071
        "--------", -- 0x3072
        "--------", -- 0x3073
        "--------", -- 0x3074
        "--------", -- 0x3075
        "--------", -- 0x3076
        "--------", -- 0x3077
        "--------", -- 0x3078
        "--------", -- 0x3079
        "--------", -- 0x307A
        "--------", -- 0x307B
        "--------", -- 0x307C
        "--------", -- 0x307D
        "--------", -- 0x307E
        "--------", -- 0x307F
        "--------", -- 0x3080
        "--------", -- 0x3081
        "--------", -- 0x3082
        "--------", -- 0x3083
        "--------", -- 0x3084
        "--------", -- 0x3085
        "--------", -- 0x3086
        "--------", -- 0x3087
        "--------", -- 0x3088
        "--------", -- 0x3089
        "--------", -- 0x308A
        "--------", -- 0x308B
        "--------", -- 0x308C
        "--------", -- 0x308D
        "--------", -- 0x308E
        "--------", -- 0x308F
        "--------", -- 0x3090
        "--------", -- 0x3091
        "--------", -- 0x3092
        "--------", -- 0x3093
        "--------", -- 0x3094
        "--------", -- 0x3095
        "--------", -- 0x3096
        "--------", -- 0x3097
        "--------", -- 0x3098
        "--------", -- 0x3099
        "--------", -- 0x309A
        "--------", -- 0x309B
        "--------", -- 0x309C
        "--------", -- 0x309D
        "--------", -- 0x309E
        "--------", -- 0x309F
        "--------", -- 0x30A0
        "--------", -- 0x30A1
        "--------", -- 0x30A2
        "--------", -- 0x30A3
        "--------", -- 0x30A4
        "--------", -- 0x30A5
        "--------", -- 0x30A6
        "--------", -- 0x30A7
        "--------", -- 0x30A8
        "--------", -- 0x30A9
        "--------", -- 0x30AA
        "--------", -- 0x30AB
        "--------", -- 0x30AC
        "--------", -- 0x30AD
        "--------", -- 0x30AE
        "--------", -- 0x30AF
        "--------", -- 0x30B0
        "--------", -- 0x30B1
        "--------", -- 0x30B2
        "--------", -- 0x30B3
        "--------", -- 0x30B4
        "--------", -- 0x30B5
        "--------", -- 0x30B6
        "--------", -- 0x30B7
        "--------", -- 0x30B8
        "--------", -- 0x30B9
        "--------", -- 0x30BA
        "--------", -- 0x30BB
        "--------", -- 0x30BC
        "--------", -- 0x30BD
        "--------", -- 0x30BE
        "--------", -- 0x30BF
        "--------", -- 0x30C0
        "--------", -- 0x30C1
        "--------", -- 0x30C2
        "--------", -- 0x30C3
        "--------", -- 0x30C4
        "--------", -- 0x30C5
        "--------", -- 0x30C6
        "--------", -- 0x30C7
        "--------", -- 0x30C8
        "--------", -- 0x30C9
        "--------", -- 0x30CA
        "--------", -- 0x30CB
        "--------", -- 0x30CC
        "--------", -- 0x30CD
        "--------", -- 0x30CE
        "--------", -- 0x30CF
        "--------", -- 0x30D0
        "--------", -- 0x30D1
        "--------", -- 0x30D2
        "--------", -- 0x30D3
        "--------", -- 0x30D4
        "--------", -- 0x30D5
        "--------", -- 0x30D6
        "--------", -- 0x30D7
        "--------", -- 0x30D8
        "--------", -- 0x30D9
        "--------", -- 0x30DA
        "--------", -- 0x30DB
        "--------", -- 0x30DC
        "--------", -- 0x30DD
        "--------", -- 0x30DE
        "--------", -- 0x30DF
        "--------", -- 0x30E0
        "--------", -- 0x30E1
        "--------", -- 0x30E2
        "--------", -- 0x30E3
        "--------", -- 0x30E4
        "--------", -- 0x30E5
        "--------", -- 0x30E6
        "--------", -- 0x30E7
        "--------", -- 0x30E8
        "--------", -- 0x30E9
        "--------", -- 0x30EA
        "--------", -- 0x30EB
        "--------", -- 0x30EC
        "--------", -- 0x30ED
        "--------", -- 0x30EE
        "--------", -- 0x30EF
        "--------", -- 0x30F0
        "--------", -- 0x30F1
        "--------", -- 0x30F2
        "--------", -- 0x30F3
        "--------", -- 0x30F4
        "--------", -- 0x30F5
        "--------", -- 0x30F6
        "--------", -- 0x30F7
        "--------", -- 0x30F8
        "--------", -- 0x30F9
        "--------", -- 0x30FA
        "--------", -- 0x30FB
        "--------", -- 0x30FC
        "--------", -- 0x30FD
        "--------", -- 0x30FE
        "--------", -- 0x30FF
        "--------", -- 0x3100
        "--------", -- 0x3101
        "--------", -- 0x3102
        "--------", -- 0x3103
        "--------", -- 0x3104
        "--------", -- 0x3105
        "--------", -- 0x3106
        "--------", -- 0x3107
        "--------", -- 0x3108
        "--------", -- 0x3109
        "--------", -- 0x310A
        "--------", -- 0x310B
        "--------", -- 0x310C
        "--------", -- 0x310D
        "--------", -- 0x310E
        "--------", -- 0x310F
        "--------", -- 0x3110
        "--------", -- 0x3111
        "--------", -- 0x3112
        "--------", -- 0x3113
        "--------", -- 0x3114
        "--------", -- 0x3115
        "--------", -- 0x3116
        "--------", -- 0x3117
        "--------", -- 0x3118
        "--------", -- 0x3119
        "--------", -- 0x311A
        "--------", -- 0x311B
        "--------", -- 0x311C
        "--------", -- 0x311D
        "--------", -- 0x311E
        "--------", -- 0x311F
        "--------", -- 0x3120
        "--------", -- 0x3121
        "--------", -- 0x3122
        "--------", -- 0x3123
        "--------", -- 0x3124
        "--------", -- 0x3125
        "--------", -- 0x3126
        "--------", -- 0x3127
        "--------", -- 0x3128
        "--------", -- 0x3129
        "--------", -- 0x312A
        "--------", -- 0x312B
        "--------", -- 0x312C
        "--------", -- 0x312D
        "--------", -- 0x312E
        "--------", -- 0x312F
        "--------", -- 0x3130
        "--------", -- 0x3131
        "--------", -- 0x3132
        "--------", -- 0x3133
        "--------", -- 0x3134
        "--------", -- 0x3135
        "--------", -- 0x3136
        "--------", -- 0x3137
        "--------", -- 0x3138
        "--------", -- 0x3139
        "--------", -- 0x313A
        "--------", -- 0x313B
        "--------", -- 0x313C
        "--------", -- 0x313D
        "--------", -- 0x313E
        "--------", -- 0x313F
        "--------", -- 0x3140
        "--------", -- 0x3141
        "--------", -- 0x3142
        "--------", -- 0x3143
        "--------", -- 0x3144
        "--------", -- 0x3145
        "--------", -- 0x3146
        "--------", -- 0x3147
        "--------", -- 0x3148
        "--------", -- 0x3149
        "--------", -- 0x314A
        "--------", -- 0x314B
        "--------", -- 0x314C
        "--------", -- 0x314D
        "--------", -- 0x314E
        "--------", -- 0x314F
        "--------", -- 0x3150
        "--------", -- 0x3151
        "--------", -- 0x3152
        "--------", -- 0x3153
        "--------", -- 0x3154
        "--------", -- 0x3155
        "--------", -- 0x3156
        "--------", -- 0x3157
        "--------", -- 0x3158
        "--------", -- 0x3159
        "--------", -- 0x315A
        "--------", -- 0x315B
        "--------", -- 0x315C
        "--------", -- 0x315D
        "--------", -- 0x315E
        "--------", -- 0x315F
        "--------", -- 0x3160
        "--------", -- 0x3161
        "--------", -- 0x3162
        "--------", -- 0x3163
        "--------", -- 0x3164
        "--------", -- 0x3165
        "--------", -- 0x3166
        "--------", -- 0x3167
        "--------", -- 0x3168
        "--------", -- 0x3169
        "--------", -- 0x316A
        "--------", -- 0x316B
        "--------", -- 0x316C
        "--------", -- 0x316D
        "--------", -- 0x316E
        "--------", -- 0x316F
        "--------", -- 0x3170
        "--------", -- 0x3171
        "--------", -- 0x3172
        "--------", -- 0x3173
        "--------", -- 0x3174
        "--------", -- 0x3175
        "--------", -- 0x3176
        "--------", -- 0x3177
        "--------", -- 0x3178
        "--------", -- 0x3179
        "--------", -- 0x317A
        "--------", -- 0x317B
        "--------", -- 0x317C
        "--------", -- 0x317D
        "--------", -- 0x317E
        "--------", -- 0x317F
        "--------", -- 0x3180
        "--------", -- 0x3181
        "--------", -- 0x3182
        "--------", -- 0x3183
        "--------", -- 0x3184
        "--------", -- 0x3185
        "--------", -- 0x3186
        "--------", -- 0x3187
        "--------", -- 0x3188
        "--------", -- 0x3189
        "--------", -- 0x318A
        "--------", -- 0x318B
        "--------", -- 0x318C
        "--------", -- 0x318D
        "--------", -- 0x318E
        "--------", -- 0x318F
        "--------", -- 0x3190
        "--------", -- 0x3191
        "--------", -- 0x3192
        "--------", -- 0x3193
        "--------", -- 0x3194
        "--------", -- 0x3195
        "--------", -- 0x3196
        "--------", -- 0x3197
        "--------", -- 0x3198
        "--------", -- 0x3199
        "--------", -- 0x319A
        "--------", -- 0x319B
        "--------", -- 0x319C
        "--------", -- 0x319D
        "--------", -- 0x319E
        "--------", -- 0x319F
        "--------", -- 0x31A0
        "--------", -- 0x31A1
        "--------", -- 0x31A2
        "--------", -- 0x31A3
        "--------", -- 0x31A4
        "--------", -- 0x31A5
        "--------", -- 0x31A6
        "--------", -- 0x31A7
        "--------", -- 0x31A8
        "--------", -- 0x31A9
        "--------", -- 0x31AA
        "--------", -- 0x31AB
        "--------", -- 0x31AC
        "--------", -- 0x31AD
        "--------", -- 0x31AE
        "--------", -- 0x31AF
        "--------", -- 0x31B0
        "--------", -- 0x31B1
        "--------", -- 0x31B2
        "--------", -- 0x31B3
        "--------", -- 0x31B4
        "--------", -- 0x31B5
        "--------", -- 0x31B6
        "--------", -- 0x31B7
        "--------", -- 0x31B8
        "--------", -- 0x31B9
        "--------", -- 0x31BA
        "--------", -- 0x31BB
        "--------", -- 0x31BC
        "--------", -- 0x31BD
        "--------", -- 0x31BE
        "--------", -- 0x31BF
        "--------", -- 0x31C0
        "--------", -- 0x31C1
        "--------", -- 0x31C2
        "--------", -- 0x31C3
        "--------", -- 0x31C4
        "--------", -- 0x31C5
        "--------", -- 0x31C6
        "--------", -- 0x31C7
        "--------", -- 0x31C8
        "--------", -- 0x31C9
        "--------", -- 0x31CA
        "--------", -- 0x31CB
        "--------", -- 0x31CC
        "--------", -- 0x31CD
        "--------", -- 0x31CE
        "--------", -- 0x31CF
        "--------", -- 0x31D0
        "--------", -- 0x31D1
        "--------", -- 0x31D2
        "--------", -- 0x31D3
        "--------", -- 0x31D4
        "--------", -- 0x31D5
        "--------", -- 0x31D6
        "--------", -- 0x31D7
        "--------", -- 0x31D8
        "--------", -- 0x31D9
        "--------", -- 0x31DA
        "--------", -- 0x31DB
        "--------", -- 0x31DC
        "--------", -- 0x31DD
        "--------", -- 0x31DE
        "--------", -- 0x31DF
        "--------", -- 0x31E0
        "--------", -- 0x31E1
        "--------", -- 0x31E2
        "--------", -- 0x31E3
        "--------", -- 0x31E4
        "--------", -- 0x31E5
        "--------", -- 0x31E6
        "--------", -- 0x31E7
        "--------", -- 0x31E8
        "--------", -- 0x31E9
        "--------", -- 0x31EA
        "--------", -- 0x31EB
        "--------", -- 0x31EC
        "--------", -- 0x31ED
        "--------", -- 0x31EE
        "--------", -- 0x31EF
        "--------", -- 0x31F0
        "--------", -- 0x31F1
        "--------", -- 0x31F2
        "--------", -- 0x31F3
        "--------", -- 0x31F4
        "--------", -- 0x31F5
        "--------", -- 0x31F6
        "--------", -- 0x31F7
        "--------", -- 0x31F8
        "--------", -- 0x31F9
        "--------", -- 0x31FA
        "--------", -- 0x31FB
        "--------", -- 0x31FC
        "--------", -- 0x31FD
        "--------", -- 0x31FE
        "--------", -- 0x31FF
        "--------", -- 0x3200
        "--------", -- 0x3201
        "--------", -- 0x3202
        "--------", -- 0x3203
        "--------", -- 0x3204
        "--------", -- 0x3205
        "--------", -- 0x3206
        "--------", -- 0x3207
        "--------", -- 0x3208
        "--------", -- 0x3209
        "--------", -- 0x320A
        "--------", -- 0x320B
        "--------", -- 0x320C
        "--------", -- 0x320D
        "--------", -- 0x320E
        "--------", -- 0x320F
        "--------", -- 0x3210
        "--------", -- 0x3211
        "--------", -- 0x3212
        "--------", -- 0x3213
        "--------", -- 0x3214
        "--------", -- 0x3215
        "--------", -- 0x3216
        "--------", -- 0x3217
        "--------", -- 0x3218
        "--------", -- 0x3219
        "--------", -- 0x321A
        "--------", -- 0x321B
        "--------", -- 0x321C
        "--------", -- 0x321D
        "--------", -- 0x321E
        "--------", -- 0x321F
        "--------", -- 0x3220
        "--------", -- 0x3221
        "--------", -- 0x3222
        "--------", -- 0x3223
        "--------", -- 0x3224
        "--------", -- 0x3225
        "--------", -- 0x3226
        "--------", -- 0x3227
        "--------", -- 0x3228
        "--------", -- 0x3229
        "--------", -- 0x322A
        "--------", -- 0x322B
        "--------", -- 0x322C
        "--------", -- 0x322D
        "--------", -- 0x322E
        "--------", -- 0x322F
        "--------", -- 0x3230
        "--------", -- 0x3231
        "--------", -- 0x3232
        "--------", -- 0x3233
        "--------", -- 0x3234
        "--------", -- 0x3235
        "--------", -- 0x3236
        "--------", -- 0x3237
        "--------", -- 0x3238
        "--------", -- 0x3239
        "--------", -- 0x323A
        "--------", -- 0x323B
        "--------", -- 0x323C
        "--------", -- 0x323D
        "--------", -- 0x323E
        "--------", -- 0x323F
        "--------", -- 0x3240
        "--------", -- 0x3241
        "--------", -- 0x3242
        "--------", -- 0x3243
        "--------", -- 0x3244
        "--------", -- 0x3245
        "--------", -- 0x3246
        "--------", -- 0x3247
        "--------", -- 0x3248
        "--------", -- 0x3249
        "--------", -- 0x324A
        "--------", -- 0x324B
        "--------", -- 0x324C
        "--------", -- 0x324D
        "--------", -- 0x324E
        "--------", -- 0x324F
        "--------", -- 0x3250
        "--------", -- 0x3251
        "--------", -- 0x3252
        "--------", -- 0x3253
        "--------", -- 0x3254
        "--------", -- 0x3255
        "--------", -- 0x3256
        "--------", -- 0x3257
        "--------", -- 0x3258
        "--------", -- 0x3259
        "--------", -- 0x325A
        "--------", -- 0x325B
        "--------", -- 0x325C
        "--------", -- 0x325D
        "--------", -- 0x325E
        "--------", -- 0x325F
        "--------", -- 0x3260
        "--------", -- 0x3261
        "--------", -- 0x3262
        "--------", -- 0x3263
        "--------", -- 0x3264
        "--------", -- 0x3265
        "--------", -- 0x3266
        "--------", -- 0x3267
        "--------", -- 0x3268
        "--------", -- 0x3269
        "--------", -- 0x326A
        "--------", -- 0x326B
        "--------", -- 0x326C
        "--------", -- 0x326D
        "--------", -- 0x326E
        "--------", -- 0x326F
        "--------", -- 0x3270
        "--------", -- 0x3271
        "--------", -- 0x3272
        "--------", -- 0x3273
        "--------", -- 0x3274
        "--------", -- 0x3275
        "--------", -- 0x3276
        "--------", -- 0x3277
        "--------", -- 0x3278
        "--------", -- 0x3279
        "--------", -- 0x327A
        "--------", -- 0x327B
        "--------", -- 0x327C
        "--------", -- 0x327D
        "--------", -- 0x327E
        "--------", -- 0x327F
        "--------", -- 0x3280
        "--------", -- 0x3281
        "--------", -- 0x3282
        "--------", -- 0x3283
        "--------", -- 0x3284
        "--------", -- 0x3285
        "--------", -- 0x3286
        "--------", -- 0x3287
        "--------", -- 0x3288
        "--------", -- 0x3289
        "--------", -- 0x328A
        "--------", -- 0x328B
        "--------", -- 0x328C
        "--------", -- 0x328D
        "--------", -- 0x328E
        "--------", -- 0x328F
        "--------", -- 0x3290
        "--------", -- 0x3291
        "--------", -- 0x3292
        "--------", -- 0x3293
        "--------", -- 0x3294
        "--------", -- 0x3295
        "--------", -- 0x3296
        "--------", -- 0x3297
        "--------", -- 0x3298
        "--------", -- 0x3299
        "--------", -- 0x329A
        "--------", -- 0x329B
        "--------", -- 0x329C
        "--------", -- 0x329D
        "--------", -- 0x329E
        "--------", -- 0x329F
        "--------", -- 0x32A0
        "--------", -- 0x32A1
        "--------", -- 0x32A2
        "--------", -- 0x32A3
        "--------", -- 0x32A4
        "--------", -- 0x32A5
        "--------", -- 0x32A6
        "--------", -- 0x32A7
        "--------", -- 0x32A8
        "--------", -- 0x32A9
        "--------", -- 0x32AA
        "--------", -- 0x32AB
        "--------", -- 0x32AC
        "--------", -- 0x32AD
        "--------", -- 0x32AE
        "--------", -- 0x32AF
        "--------", -- 0x32B0
        "--------", -- 0x32B1
        "--------", -- 0x32B2
        "--------", -- 0x32B3
        "--------", -- 0x32B4
        "--------", -- 0x32B5
        "--------", -- 0x32B6
        "--------", -- 0x32B7
        "--------", -- 0x32B8
        "--------", -- 0x32B9
        "--------", -- 0x32BA
        "--------", -- 0x32BB
        "--------", -- 0x32BC
        "--------", -- 0x32BD
        "--------", -- 0x32BE
        "--------", -- 0x32BF
        "--------", -- 0x32C0
        "--------", -- 0x32C1
        "--------", -- 0x32C2
        "--------", -- 0x32C3
        "--------", -- 0x32C4
        "--------", -- 0x32C5
        "--------", -- 0x32C6
        "--------", -- 0x32C7
        "--------", -- 0x32C8
        "--------", -- 0x32C9
        "--------", -- 0x32CA
        "--------", -- 0x32CB
        "--------", -- 0x32CC
        "--------", -- 0x32CD
        "--------", -- 0x32CE
        "--------", -- 0x32CF
        "--------", -- 0x32D0
        "--------", -- 0x32D1
        "--------", -- 0x32D2
        "--------", -- 0x32D3
        "--------", -- 0x32D4
        "--------", -- 0x32D5
        "--------", -- 0x32D6
        "--------", -- 0x32D7
        "--------", -- 0x32D8
        "--------", -- 0x32D9
        "--------", -- 0x32DA
        "--------", -- 0x32DB
        "--------", -- 0x32DC
        "--------", -- 0x32DD
        "--------", -- 0x32DE
        "--------", -- 0x32DF
        "--------", -- 0x32E0
        "--------", -- 0x32E1
        "--------", -- 0x32E2
        "--------", -- 0x32E3
        "--------", -- 0x32E4
        "--------", -- 0x32E5
        "--------", -- 0x32E6
        "--------", -- 0x32E7
        "--------", -- 0x32E8
        "--------", -- 0x32E9
        "--------", -- 0x32EA
        "--------", -- 0x32EB
        "--------", -- 0x32EC
        "--------", -- 0x32ED
        "--------", -- 0x32EE
        "--------", -- 0x32EF
        "--------", -- 0x32F0
        "--------", -- 0x32F1
        "--------", -- 0x32F2
        "--------", -- 0x32F3
        "--------", -- 0x32F4
        "--------", -- 0x32F5
        "--------", -- 0x32F6
        "--------", -- 0x32F7
        "--------", -- 0x32F8
        "--------", -- 0x32F9
        "--------", -- 0x32FA
        "--------", -- 0x32FB
        "--------", -- 0x32FC
        "--------", -- 0x32FD
        "--------", -- 0x32FE
        "--------", -- 0x32FF
        "--------", -- 0x3300
        "--------", -- 0x3301
        "--------", -- 0x3302
        "--------", -- 0x3303
        "--------", -- 0x3304
        "--------", -- 0x3305
        "--------", -- 0x3306
        "--------", -- 0x3307
        "--------", -- 0x3308
        "--------", -- 0x3309
        "--------", -- 0x330A
        "--------", -- 0x330B
        "--------", -- 0x330C
        "--------", -- 0x330D
        "--------", -- 0x330E
        "--------", -- 0x330F
        "--------", -- 0x3310
        "--------", -- 0x3311
        "--------", -- 0x3312
        "--------", -- 0x3313
        "--------", -- 0x3314
        "--------", -- 0x3315
        "--------", -- 0x3316
        "--------", -- 0x3317
        "--------", -- 0x3318
        "--------", -- 0x3319
        "--------", -- 0x331A
        "--------", -- 0x331B
        "--------", -- 0x331C
        "--------", -- 0x331D
        "--------", -- 0x331E
        "--------", -- 0x331F
        "--------", -- 0x3320
        "--------", -- 0x3321
        "--------", -- 0x3322
        "--------", -- 0x3323
        "--------", -- 0x3324
        "--------", -- 0x3325
        "--------", -- 0x3326
        "--------", -- 0x3327
        "--------", -- 0x3328
        "--------", -- 0x3329
        "--------", -- 0x332A
        "--------", -- 0x332B
        "--------", -- 0x332C
        "--------", -- 0x332D
        "--------", -- 0x332E
        "--------", -- 0x332F
        "--------", -- 0x3330
        "--------", -- 0x3331
        "--------", -- 0x3332
        "--------", -- 0x3333
        "--------", -- 0x3334
        "--------", -- 0x3335
        "--------", -- 0x3336
        "--------", -- 0x3337
        "--------", -- 0x3338
        "--------", -- 0x3339
        "--------", -- 0x333A
        "--------", -- 0x333B
        "--------", -- 0x333C
        "--------", -- 0x333D
        "--------", -- 0x333E
        "--------", -- 0x333F
        "--------", -- 0x3340
        "--------", -- 0x3341
        "--------", -- 0x3342
        "--------", -- 0x3343
        "--------", -- 0x3344
        "--------", -- 0x3345
        "--------", -- 0x3346
        "--------", -- 0x3347
        "--------", -- 0x3348
        "--------", -- 0x3349
        "--------", -- 0x334A
        "--------", -- 0x334B
        "--------", -- 0x334C
        "--------", -- 0x334D
        "--------", -- 0x334E
        "--------", -- 0x334F
        "--------", -- 0x3350
        "--------", -- 0x3351
        "--------", -- 0x3352
        "--------", -- 0x3353
        "--------", -- 0x3354
        "--------", -- 0x3355
        "--------", -- 0x3356
        "--------", -- 0x3357
        "--------", -- 0x3358
        "--------", -- 0x3359
        "--------", -- 0x335A
        "--------", -- 0x335B
        "--------", -- 0x335C
        "--------", -- 0x335D
        "--------", -- 0x335E
        "--------", -- 0x335F
        "--------", -- 0x3360
        "--------", -- 0x3361
        "--------", -- 0x3362
        "--------", -- 0x3363
        "--------", -- 0x3364
        "--------", -- 0x3365
        "--------", -- 0x3366
        "--------", -- 0x3367
        "--------", -- 0x3368
        "--------", -- 0x3369
        "--------", -- 0x336A
        "--------", -- 0x336B
        "--------", -- 0x336C
        "--------", -- 0x336D
        "--------", -- 0x336E
        "--------", -- 0x336F
        "--------", -- 0x3370
        "--------", -- 0x3371
        "--------", -- 0x3372
        "--------", -- 0x3373
        "--------", -- 0x3374
        "--------", -- 0x3375
        "--------", -- 0x3376
        "--------", -- 0x3377
        "--------", -- 0x3378
        "--------", -- 0x3379
        "--------", -- 0x337A
        "--------", -- 0x337B
        "--------", -- 0x337C
        "--------", -- 0x337D
        "--------", -- 0x337E
        "--------", -- 0x337F
        "--------", -- 0x3380
        "--------", -- 0x3381
        "--------", -- 0x3382
        "--------", -- 0x3383
        "--------", -- 0x3384
        "--------", -- 0x3385
        "--------", -- 0x3386
        "--------", -- 0x3387
        "--------", -- 0x3388
        "--------", -- 0x3389
        "--------", -- 0x338A
        "--------", -- 0x338B
        "--------", -- 0x338C
        "--------", -- 0x338D
        "--------", -- 0x338E
        "--------", -- 0x338F
        "--------", -- 0x3390
        "--------", -- 0x3391
        "--------", -- 0x3392
        "--------", -- 0x3393
        "--------", -- 0x3394
        "--------", -- 0x3395
        "--------", -- 0x3396
        "--------", -- 0x3397
        "--------", -- 0x3398
        "--------", -- 0x3399
        "--------", -- 0x339A
        "--------", -- 0x339B
        "--------", -- 0x339C
        "--------", -- 0x339D
        "--------", -- 0x339E
        "--------", -- 0x339F
        "--------", -- 0x33A0
        "--------", -- 0x33A1
        "--------", -- 0x33A2
        "--------", -- 0x33A3
        "--------", -- 0x33A4
        "--------", -- 0x33A5
        "--------", -- 0x33A6
        "--------", -- 0x33A7
        "--------", -- 0x33A8
        "--------", -- 0x33A9
        "--------", -- 0x33AA
        "--------", -- 0x33AB
        "--------", -- 0x33AC
        "--------", -- 0x33AD
        "--------", -- 0x33AE
        "--------", -- 0x33AF
        "--------", -- 0x33B0
        "--------", -- 0x33B1
        "--------", -- 0x33B2
        "--------", -- 0x33B3
        "--------", -- 0x33B4
        "--------", -- 0x33B5
        "--------", -- 0x33B6
        "--------", -- 0x33B7
        "--------", -- 0x33B8
        "--------", -- 0x33B9
        "--------", -- 0x33BA
        "--------", -- 0x33BB
        "--------", -- 0x33BC
        "--------", -- 0x33BD
        "--------", -- 0x33BE
        "--------", -- 0x33BF
        "--------", -- 0x33C0
        "--------", -- 0x33C1
        "--------", -- 0x33C2
        "--------", -- 0x33C3
        "--------", -- 0x33C4
        "--------", -- 0x33C5
        "--------", -- 0x33C6
        "--------", -- 0x33C7
        "--------", -- 0x33C8
        "--------", -- 0x33C9
        "--------", -- 0x33CA
        "--------", -- 0x33CB
        "--------", -- 0x33CC
        "--------", -- 0x33CD
        "--------", -- 0x33CE
        "--------", -- 0x33CF
        "--------", -- 0x33D0
        "--------", -- 0x33D1
        "--------", -- 0x33D2
        "--------", -- 0x33D3
        "--------", -- 0x33D4
        "--------", -- 0x33D5
        "--------", -- 0x33D6
        "--------", -- 0x33D7
        "--------", -- 0x33D8
        "--------", -- 0x33D9
        "--------", -- 0x33DA
        "--------", -- 0x33DB
        "--------", -- 0x33DC
        "--------", -- 0x33DD
        "--------", -- 0x33DE
        "--------", -- 0x33DF
        "--------", -- 0x33E0
        "--------", -- 0x33E1
        "--------", -- 0x33E2
        "--------", -- 0x33E3
        "--------", -- 0x33E4
        "--------", -- 0x33E5
        "--------", -- 0x33E6
        "--------", -- 0x33E7
        "--------", -- 0x33E8
        "--------", -- 0x33E9
        "--------", -- 0x33EA
        "--------", -- 0x33EB
        "--------", -- 0x33EC
        "--------", -- 0x33ED
        "--------", -- 0x33EE
        "--------", -- 0x33EF
        "--------", -- 0x33F0
        "--------", -- 0x33F1
        "--------", -- 0x33F2
        "--------", -- 0x33F3
        "--------", -- 0x33F4
        "--------", -- 0x33F5
        "--------", -- 0x33F6
        "--------", -- 0x33F7
        "--------", -- 0x33F8
        "--------", -- 0x33F9
        "--------", -- 0x33FA
        "--------", -- 0x33FB
        "--------", -- 0x33FC
        "--------", -- 0x33FD
        "--------", -- 0x33FE
        "--------", -- 0x33FF
        "--------", -- 0x3400
        "--------", -- 0x3401
        "--------", -- 0x3402
        "--------", -- 0x3403
        "--------", -- 0x3404
        "--------", -- 0x3405
        "--------", -- 0x3406
        "--------", -- 0x3407
        "--------", -- 0x3408
        "--------", -- 0x3409
        "--------", -- 0x340A
        "--------", -- 0x340B
        "--------", -- 0x340C
        "--------", -- 0x340D
        "--------", -- 0x340E
        "--------", -- 0x340F
        "--------", -- 0x3410
        "--------", -- 0x3411
        "--------", -- 0x3412
        "--------", -- 0x3413
        "--------", -- 0x3414
        "--------", -- 0x3415
        "--------", -- 0x3416
        "--------", -- 0x3417
        "--------", -- 0x3418
        "--------", -- 0x3419
        "--------", -- 0x341A
        "--------", -- 0x341B
        "--------", -- 0x341C
        "--------", -- 0x341D
        "--------", -- 0x341E
        "--------", -- 0x341F
        "--------", -- 0x3420
        "--------", -- 0x3421
        "--------", -- 0x3422
        "--------", -- 0x3423
        "--------", -- 0x3424
        "--------", -- 0x3425
        "--------", -- 0x3426
        "--------", -- 0x3427
        "--------", -- 0x3428
        "--------", -- 0x3429
        "--------", -- 0x342A
        "--------", -- 0x342B
        "--------", -- 0x342C
        "--------", -- 0x342D
        "--------", -- 0x342E
        "--------", -- 0x342F
        "--------", -- 0x3430
        "--------", -- 0x3431
        "--------", -- 0x3432
        "--------", -- 0x3433
        "--------", -- 0x3434
        "--------", -- 0x3435
        "--------", -- 0x3436
        "--------", -- 0x3437
        "--------", -- 0x3438
        "--------", -- 0x3439
        "--------", -- 0x343A
        "--------", -- 0x343B
        "--------", -- 0x343C
        "--------", -- 0x343D
        "--------", -- 0x343E
        "--------", -- 0x343F
        "--------", -- 0x3440
        "--------", -- 0x3441
        "--------", -- 0x3442
        "--------", -- 0x3443
        "--------", -- 0x3444
        "--------", -- 0x3445
        "--------", -- 0x3446
        "--------", -- 0x3447
        "--------", -- 0x3448
        "--------", -- 0x3449
        "--------", -- 0x344A
        "--------", -- 0x344B
        "--------", -- 0x344C
        "--------", -- 0x344D
        "--------", -- 0x344E
        "--------", -- 0x344F
        "--------", -- 0x3450
        "--------", -- 0x3451
        "--------", -- 0x3452
        "--------", -- 0x3453
        "--------", -- 0x3454
        "--------", -- 0x3455
        "--------", -- 0x3456
        "--------", -- 0x3457
        "--------", -- 0x3458
        "--------", -- 0x3459
        "--------", -- 0x345A
        "--------", -- 0x345B
        "--------", -- 0x345C
        "--------", -- 0x345D
        "--------", -- 0x345E
        "--------", -- 0x345F
        "--------", -- 0x3460
        "--------", -- 0x3461
        "--------", -- 0x3462
        "--------", -- 0x3463
        "--------", -- 0x3464
        "--------", -- 0x3465
        "--------", -- 0x3466
        "--------", -- 0x3467
        "--------", -- 0x3468
        "--------", -- 0x3469
        "--------", -- 0x346A
        "--------", -- 0x346B
        "--------", -- 0x346C
        "--------", -- 0x346D
        "--------", -- 0x346E
        "--------", -- 0x346F
        "--------", -- 0x3470
        "--------", -- 0x3471
        "--------", -- 0x3472
        "--------", -- 0x3473
        "--------", -- 0x3474
        "--------", -- 0x3475
        "--------", -- 0x3476
        "--------", -- 0x3477
        "--------", -- 0x3478
        "--------", -- 0x3479
        "--------", -- 0x347A
        "--------", -- 0x347B
        "--------", -- 0x347C
        "--------", -- 0x347D
        "--------", -- 0x347E
        "--------", -- 0x347F
        "--------", -- 0x3480
        "--------", -- 0x3481
        "--------", -- 0x3482
        "--------", -- 0x3483
        "--------", -- 0x3484
        "--------", -- 0x3485
        "--------", -- 0x3486
        "--------", -- 0x3487
        "--------", -- 0x3488
        "--------", -- 0x3489
        "--------", -- 0x348A
        "--------", -- 0x348B
        "--------", -- 0x348C
        "--------", -- 0x348D
        "--------", -- 0x348E
        "--------", -- 0x348F
        "--------", -- 0x3490
        "--------", -- 0x3491
        "--------", -- 0x3492
        "--------", -- 0x3493
        "--------", -- 0x3494
        "--------", -- 0x3495
        "--------", -- 0x3496
        "--------", -- 0x3497
        "--------", -- 0x3498
        "--------", -- 0x3499
        "--------", -- 0x349A
        "--------", -- 0x349B
        "--------", -- 0x349C
        "--------", -- 0x349D
        "--------", -- 0x349E
        "--------", -- 0x349F
        "--------", -- 0x34A0
        "--------", -- 0x34A1
        "--------", -- 0x34A2
        "--------", -- 0x34A3
        "--------", -- 0x34A4
        "--------", -- 0x34A5
        "--------", -- 0x34A6
        "--------", -- 0x34A7
        "--------", -- 0x34A8
        "--------", -- 0x34A9
        "--------", -- 0x34AA
        "--------", -- 0x34AB
        "--------", -- 0x34AC
        "--------", -- 0x34AD
        "--------", -- 0x34AE
        "--------", -- 0x34AF
        "--------", -- 0x34B0
        "--------", -- 0x34B1
        "--------", -- 0x34B2
        "--------", -- 0x34B3
        "--------", -- 0x34B4
        "--------", -- 0x34B5
        "--------", -- 0x34B6
        "--------", -- 0x34B7
        "--------", -- 0x34B8
        "--------", -- 0x34B9
        "--------", -- 0x34BA
        "--------", -- 0x34BB
        "--------", -- 0x34BC
        "--------", -- 0x34BD
        "--------", -- 0x34BE
        "--------", -- 0x34BF
        "--------", -- 0x34C0
        "--------", -- 0x34C1
        "--------", -- 0x34C2
        "--------", -- 0x34C3
        "--------", -- 0x34C4
        "--------", -- 0x34C5
        "--------", -- 0x34C6
        "--------", -- 0x34C7
        "--------", -- 0x34C8
        "--------", -- 0x34C9
        "--------", -- 0x34CA
        "--------", -- 0x34CB
        "--------", -- 0x34CC
        "--------", -- 0x34CD
        "--------", -- 0x34CE
        "--------", -- 0x34CF
        "--------", -- 0x34D0
        "--------", -- 0x34D1
        "--------", -- 0x34D2
        "--------", -- 0x34D3
        "--------", -- 0x34D4
        "--------", -- 0x34D5
        "--------", -- 0x34D6
        "--------", -- 0x34D7
        "--------", -- 0x34D8
        "--------", -- 0x34D9
        "--------", -- 0x34DA
        "--------", -- 0x34DB
        "--------", -- 0x34DC
        "--------", -- 0x34DD
        "--------", -- 0x34DE
        "--------", -- 0x34DF
        "--------", -- 0x34E0
        "--------", -- 0x34E1
        "--------", -- 0x34E2
        "--------", -- 0x34E3
        "--------", -- 0x34E4
        "--------", -- 0x34E5
        "--------", -- 0x34E6
        "--------", -- 0x34E7
        "--------", -- 0x34E8
        "--------", -- 0x34E9
        "--------", -- 0x34EA
        "--------", -- 0x34EB
        "--------", -- 0x34EC
        "--------", -- 0x34ED
        "--------", -- 0x34EE
        "--------", -- 0x34EF
        "--------", -- 0x34F0
        "--------", -- 0x34F1
        "--------", -- 0x34F2
        "--------", -- 0x34F3
        "--------", -- 0x34F4
        "--------", -- 0x34F5
        "--------", -- 0x34F6
        "--------", -- 0x34F7
        "--------", -- 0x34F8
        "--------", -- 0x34F9
        "--------", -- 0x34FA
        "--------", -- 0x34FB
        "--------", -- 0x34FC
        "--------", -- 0x34FD
        "--------", -- 0x34FE
        "--------", -- 0x34FF
        "--------", -- 0x3500
        "--------", -- 0x3501
        "--------", -- 0x3502
        "--------", -- 0x3503
        "--------", -- 0x3504
        "--------", -- 0x3505
        "--------", -- 0x3506
        "--------", -- 0x3507
        "--------", -- 0x3508
        "--------", -- 0x3509
        "--------", -- 0x350A
        "--------", -- 0x350B
        "--------", -- 0x350C
        "--------", -- 0x350D
        "--------", -- 0x350E
        "--------", -- 0x350F
        "--------", -- 0x3510
        "--------", -- 0x3511
        "--------", -- 0x3512
        "--------", -- 0x3513
        "--------", -- 0x3514
        "--------", -- 0x3515
        "--------", -- 0x3516
        "--------", -- 0x3517
        "--------", -- 0x3518
        "--------", -- 0x3519
        "--------", -- 0x351A
        "--------", -- 0x351B
        "--------", -- 0x351C
        "--------", -- 0x351D
        "--------", -- 0x351E
        "--------", -- 0x351F
        "--------", -- 0x3520
        "--------", -- 0x3521
        "--------", -- 0x3522
        "--------", -- 0x3523
        "--------", -- 0x3524
        "--------", -- 0x3525
        "--------", -- 0x3526
        "--------", -- 0x3527
        "--------", -- 0x3528
        "--------", -- 0x3529
        "--------", -- 0x352A
        "--------", -- 0x352B
        "--------", -- 0x352C
        "--------", -- 0x352D
        "--------", -- 0x352E
        "--------", -- 0x352F
        "--------", -- 0x3530
        "--------", -- 0x3531
        "--------", -- 0x3532
        "--------", -- 0x3533
        "--------", -- 0x3534
        "--------", -- 0x3535
        "--------", -- 0x3536
        "--------", -- 0x3537
        "--------", -- 0x3538
        "--------", -- 0x3539
        "--------", -- 0x353A
        "--------", -- 0x353B
        "--------", -- 0x353C
        "--------", -- 0x353D
        "--------", -- 0x353E
        "--------", -- 0x353F
        "--------", -- 0x3540
        "--------", -- 0x3541
        "--------", -- 0x3542
        "--------", -- 0x3543
        "--------", -- 0x3544
        "--------", -- 0x3545
        "--------", -- 0x3546
        "--------", -- 0x3547
        "--------", -- 0x3548
        "--------", -- 0x3549
        "--------", -- 0x354A
        "--------", -- 0x354B
        "--------", -- 0x354C
        "--------", -- 0x354D
        "--------", -- 0x354E
        "--------", -- 0x354F
        "--------", -- 0x3550
        "--------", -- 0x3551
        "--------", -- 0x3552
        "--------", -- 0x3553
        "--------", -- 0x3554
        "--------", -- 0x3555
        "--------", -- 0x3556
        "--------", -- 0x3557
        "--------", -- 0x3558
        "--------", -- 0x3559
        "--------", -- 0x355A
        "--------", -- 0x355B
        "--------", -- 0x355C
        "--------", -- 0x355D
        "--------", -- 0x355E
        "--------", -- 0x355F
        "--------", -- 0x3560
        "--------", -- 0x3561
        "--------", -- 0x3562
        "--------", -- 0x3563
        "--------", -- 0x3564
        "--------", -- 0x3565
        "--------", -- 0x3566
        "--------", -- 0x3567
        "--------", -- 0x3568
        "--------", -- 0x3569
        "--------", -- 0x356A
        "--------", -- 0x356B
        "--------", -- 0x356C
        "--------", -- 0x356D
        "--------", -- 0x356E
        "--------", -- 0x356F
        "--------", -- 0x3570
        "--------", -- 0x3571
        "--------", -- 0x3572
        "--------", -- 0x3573
        "--------", -- 0x3574
        "--------", -- 0x3575
        "--------", -- 0x3576
        "--------", -- 0x3577
        "--------", -- 0x3578
        "--------", -- 0x3579
        "--------", -- 0x357A
        "--------", -- 0x357B
        "--------", -- 0x357C
        "--------", -- 0x357D
        "--------", -- 0x357E
        "--------", -- 0x357F
        "--------", -- 0x3580
        "--------", -- 0x3581
        "--------", -- 0x3582
        "--------", -- 0x3583
        "--------", -- 0x3584
        "--------", -- 0x3585
        "--------", -- 0x3586
        "--------", -- 0x3587
        "--------", -- 0x3588
        "--------", -- 0x3589
        "--------", -- 0x358A
        "--------", -- 0x358B
        "--------", -- 0x358C
        "--------", -- 0x358D
        "--------", -- 0x358E
        "--------", -- 0x358F
        "--------", -- 0x3590
        "--------", -- 0x3591
        "--------", -- 0x3592
        "--------", -- 0x3593
        "--------", -- 0x3594
        "--------", -- 0x3595
        "--------", -- 0x3596
        "--------", -- 0x3597
        "--------", -- 0x3598
        "--------", -- 0x3599
        "--------", -- 0x359A
        "--------", -- 0x359B
        "--------", -- 0x359C
        "--------", -- 0x359D
        "--------", -- 0x359E
        "--------", -- 0x359F
        "--------", -- 0x35A0
        "--------", -- 0x35A1
        "--------", -- 0x35A2
        "--------", -- 0x35A3
        "--------", -- 0x35A4
        "--------", -- 0x35A5
        "--------", -- 0x35A6
        "--------", -- 0x35A7
        "--------", -- 0x35A8
        "--------", -- 0x35A9
        "--------", -- 0x35AA
        "--------", -- 0x35AB
        "--------", -- 0x35AC
        "--------", -- 0x35AD
        "--------", -- 0x35AE
        "--------", -- 0x35AF
        "--------", -- 0x35B0
        "--------", -- 0x35B1
        "--------", -- 0x35B2
        "--------", -- 0x35B3
        "--------", -- 0x35B4
        "--------", -- 0x35B5
        "--------", -- 0x35B6
        "--------", -- 0x35B7
        "--------", -- 0x35B8
        "--------", -- 0x35B9
        "--------", -- 0x35BA
        "--------", -- 0x35BB
        "--------", -- 0x35BC
        "--------", -- 0x35BD
        "--------", -- 0x35BE
        "--------", -- 0x35BF
        "--------", -- 0x35C0
        "--------", -- 0x35C1
        "--------", -- 0x35C2
        "--------", -- 0x35C3
        "--------", -- 0x35C4
        "--------", -- 0x35C5
        "--------", -- 0x35C6
        "--------", -- 0x35C7
        "--------", -- 0x35C8
        "--------", -- 0x35C9
        "--------", -- 0x35CA
        "--------", -- 0x35CB
        "--------", -- 0x35CC
        "--------", -- 0x35CD
        "--------", -- 0x35CE
        "--------", -- 0x35CF
        "--------", -- 0x35D0
        "--------", -- 0x35D1
        "--------", -- 0x35D2
        "--------", -- 0x35D3
        "--------", -- 0x35D4
        "--------", -- 0x35D5
        "--------", -- 0x35D6
        "--------", -- 0x35D7
        "--------", -- 0x35D8
        "--------", -- 0x35D9
        "--------", -- 0x35DA
        "--------", -- 0x35DB
        "--------", -- 0x35DC
        "--------", -- 0x35DD
        "--------", -- 0x35DE
        "--------", -- 0x35DF
        "--------", -- 0x35E0
        "--------", -- 0x35E1
        "--------", -- 0x35E2
        "--------", -- 0x35E3
        "--------", -- 0x35E4
        "--------", -- 0x35E5
        "--------", -- 0x35E6
        "--------", -- 0x35E7
        "--------", -- 0x35E8
        "--------", -- 0x35E9
        "--------", -- 0x35EA
        "--------", -- 0x35EB
        "--------", -- 0x35EC
        "--------", -- 0x35ED
        "--------", -- 0x35EE
        "--------", -- 0x35EF
        "--------", -- 0x35F0
        "--------", -- 0x35F1
        "--------", -- 0x35F2
        "--------", -- 0x35F3
        "--------", -- 0x35F4
        "--------", -- 0x35F5
        "--------", -- 0x35F6
        "--------", -- 0x35F7
        "--------", -- 0x35F8
        "--------", -- 0x35F9
        "--------", -- 0x35FA
        "--------", -- 0x35FB
        "--------", -- 0x35FC
        "--------", -- 0x35FD
        "--------", -- 0x35FE
        "--------", -- 0x35FF
        "--------", -- 0x3600
        "--------", -- 0x3601
        "--------", -- 0x3602
        "--------", -- 0x3603
        "--------", -- 0x3604
        "--------", -- 0x3605
        "--------", -- 0x3606
        "--------", -- 0x3607
        "--------", -- 0x3608
        "--------", -- 0x3609
        "--------", -- 0x360A
        "--------", -- 0x360B
        "--------", -- 0x360C
        "--------", -- 0x360D
        "--------", -- 0x360E
        "--------", -- 0x360F
        "--------", -- 0x3610
        "--------", -- 0x3611
        "--------", -- 0x3612
        "--------", -- 0x3613
        "--------", -- 0x3614
        "--------", -- 0x3615
        "--------", -- 0x3616
        "--------", -- 0x3617
        "--------", -- 0x3618
        "--------", -- 0x3619
        "--------", -- 0x361A
        "--------", -- 0x361B
        "--------", -- 0x361C
        "--------", -- 0x361D
        "--------", -- 0x361E
        "--------", -- 0x361F
        "--------", -- 0x3620
        "--------", -- 0x3621
        "--------", -- 0x3622
        "--------", -- 0x3623
        "--------", -- 0x3624
        "--------", -- 0x3625
        "--------", -- 0x3626
        "--------", -- 0x3627
        "--------", -- 0x3628
        "--------", -- 0x3629
        "--------", -- 0x362A
        "--------", -- 0x362B
        "--------", -- 0x362C
        "--------", -- 0x362D
        "--------", -- 0x362E
        "--------", -- 0x362F
        "--------", -- 0x3630
        "--------", -- 0x3631
        "--------", -- 0x3632
        "--------", -- 0x3633
        "--------", -- 0x3634
        "--------", -- 0x3635
        "--------", -- 0x3636
        "--------", -- 0x3637
        "--------", -- 0x3638
        "--------", -- 0x3639
        "--------", -- 0x363A
        "--------", -- 0x363B
        "--------", -- 0x363C
        "--------", -- 0x363D
        "--------", -- 0x363E
        "--------", -- 0x363F
        "--------", -- 0x3640
        "--------", -- 0x3641
        "--------", -- 0x3642
        "--------", -- 0x3643
        "--------", -- 0x3644
        "--------", -- 0x3645
        "--------", -- 0x3646
        "--------", -- 0x3647
        "--------", -- 0x3648
        "--------", -- 0x3649
        "--------", -- 0x364A
        "--------", -- 0x364B
        "--------", -- 0x364C
        "--------", -- 0x364D
        "--------", -- 0x364E
        "--------", -- 0x364F
        "--------", -- 0x3650
        "--------", -- 0x3651
        "--------", -- 0x3652
        "--------", -- 0x3653
        "--------", -- 0x3654
        "--------", -- 0x3655
        "--------", -- 0x3656
        "--------", -- 0x3657
        "--------", -- 0x3658
        "--------", -- 0x3659
        "--------", -- 0x365A
        "--------", -- 0x365B
        "--------", -- 0x365C
        "--------", -- 0x365D
        "--------", -- 0x365E
        "--------", -- 0x365F
        "--------", -- 0x3660
        "--------", -- 0x3661
        "--------", -- 0x3662
        "--------", -- 0x3663
        "--------", -- 0x3664
        "--------", -- 0x3665
        "--------", -- 0x3666
        "--------", -- 0x3667
        "--------", -- 0x3668
        "--------", -- 0x3669
        "--------", -- 0x366A
        "--------", -- 0x366B
        "--------", -- 0x366C
        "--------", -- 0x366D
        "--------", -- 0x366E
        "--------", -- 0x366F
        "--------", -- 0x3670
        "--------", -- 0x3671
        "--------", -- 0x3672
        "--------", -- 0x3673
        "--------", -- 0x3674
        "--------", -- 0x3675
        "--------", -- 0x3676
        "--------", -- 0x3677
        "--------", -- 0x3678
        "--------", -- 0x3679
        "--------", -- 0x367A
        "--------", -- 0x367B
        "--------", -- 0x367C
        "--------", -- 0x367D
        "--------", -- 0x367E
        "--------", -- 0x367F
        "--------", -- 0x3680
        "--------", -- 0x3681
        "--------", -- 0x3682
        "--------", -- 0x3683
        "--------", -- 0x3684
        "--------", -- 0x3685
        "--------", -- 0x3686
        "--------", -- 0x3687
        "--------", -- 0x3688
        "--------", -- 0x3689
        "--------", -- 0x368A
        "--------", -- 0x368B
        "--------", -- 0x368C
        "--------", -- 0x368D
        "--------", -- 0x368E
        "--------", -- 0x368F
        "--------", -- 0x3690
        "--------", -- 0x3691
        "--------", -- 0x3692
        "--------", -- 0x3693
        "--------", -- 0x3694
        "--------", -- 0x3695
        "--------", -- 0x3696
        "--------", -- 0x3697
        "--------", -- 0x3698
        "--------", -- 0x3699
        "--------", -- 0x369A
        "--------", -- 0x369B
        "--------", -- 0x369C
        "--------", -- 0x369D
        "--------", -- 0x369E
        "--------", -- 0x369F
        "--------", -- 0x36A0
        "--------", -- 0x36A1
        "--------", -- 0x36A2
        "--------", -- 0x36A3
        "--------", -- 0x36A4
        "--------", -- 0x36A5
        "--------", -- 0x36A6
        "--------", -- 0x36A7
        "--------", -- 0x36A8
        "--------", -- 0x36A9
        "--------", -- 0x36AA
        "--------", -- 0x36AB
        "--------", -- 0x36AC
        "--------", -- 0x36AD
        "--------", -- 0x36AE
        "--------", -- 0x36AF
        "--------", -- 0x36B0
        "--------", -- 0x36B1
        "--------", -- 0x36B2
        "--------", -- 0x36B3
        "--------", -- 0x36B4
        "--------", -- 0x36B5
        "--------", -- 0x36B6
        "--------", -- 0x36B7
        "--------", -- 0x36B8
        "--------", -- 0x36B9
        "--------", -- 0x36BA
        "--------", -- 0x36BB
        "--------", -- 0x36BC
        "--------", -- 0x36BD
        "--------", -- 0x36BE
        "--------", -- 0x36BF
        "--------", -- 0x36C0
        "--------", -- 0x36C1
        "--------", -- 0x36C2
        "--------", -- 0x36C3
        "--------", -- 0x36C4
        "--------", -- 0x36C5
        "--------", -- 0x36C6
        "--------", -- 0x36C7
        "--------", -- 0x36C8
        "--------", -- 0x36C9
        "--------", -- 0x36CA
        "--------", -- 0x36CB
        "--------", -- 0x36CC
        "--------", -- 0x36CD
        "--------", -- 0x36CE
        "--------", -- 0x36CF
        "--------", -- 0x36D0
        "--------", -- 0x36D1
        "--------", -- 0x36D2
        "--------", -- 0x36D3
        "--------", -- 0x36D4
        "--------", -- 0x36D5
        "--------", -- 0x36D6
        "--------", -- 0x36D7
        "--------", -- 0x36D8
        "--------", -- 0x36D9
        "--------", -- 0x36DA
        "--------", -- 0x36DB
        "--------", -- 0x36DC
        "--------", -- 0x36DD
        "--------", -- 0x36DE
        "--------", -- 0x36DF
        "--------", -- 0x36E0
        "--------", -- 0x36E1
        "--------", -- 0x36E2
        "--------", -- 0x36E3
        "--------", -- 0x36E4
        "--------", -- 0x36E5
        "--------", -- 0x36E6
        "--------", -- 0x36E7
        "--------", -- 0x36E8
        "--------", -- 0x36E9
        "--------", -- 0x36EA
        "--------", -- 0x36EB
        "--------", -- 0x36EC
        "--------", -- 0x36ED
        "--------", -- 0x36EE
        "--------", -- 0x36EF
        "--------", -- 0x36F0
        "--------", -- 0x36F1
        "--------", -- 0x36F2
        "--------", -- 0x36F3
        "--------", -- 0x36F4
        "--------", -- 0x36F5
        "--------", -- 0x36F6
        "--------", -- 0x36F7
        "--------", -- 0x36F8
        "--------", -- 0x36F9
        "--------", -- 0x36FA
        "--------", -- 0x36FB
        "--------", -- 0x36FC
        "--------", -- 0x36FD
        "--------", -- 0x36FE
        "--------", -- 0x36FF
        "--------", -- 0x3700
        "--------", -- 0x3701
        "--------", -- 0x3702
        "--------", -- 0x3703
        "--------", -- 0x3704
        "--------", -- 0x3705
        "--------", -- 0x3706
        "--------", -- 0x3707
        "--------", -- 0x3708
        "--------", -- 0x3709
        "--------", -- 0x370A
        "--------", -- 0x370B
        "--------", -- 0x370C
        "--------", -- 0x370D
        "--------", -- 0x370E
        "--------", -- 0x370F
        "--------", -- 0x3710
        "--------", -- 0x3711
        "--------", -- 0x3712
        "--------", -- 0x3713
        "--------", -- 0x3714
        "--------", -- 0x3715
        "--------", -- 0x3716
        "--------", -- 0x3717
        "--------", -- 0x3718
        "--------", -- 0x3719
        "--------", -- 0x371A
        "--------", -- 0x371B
        "--------", -- 0x371C
        "--------", -- 0x371D
        "--------", -- 0x371E
        "--------", -- 0x371F
        "--------", -- 0x3720
        "--------", -- 0x3721
        "--------", -- 0x3722
        "--------", -- 0x3723
        "--------", -- 0x3724
        "--------", -- 0x3725
        "--------", -- 0x3726
        "--------", -- 0x3727
        "--------", -- 0x3728
        "--------", -- 0x3729
        "--------", -- 0x372A
        "--------", -- 0x372B
        "--------", -- 0x372C
        "--------", -- 0x372D
        "--------", -- 0x372E
        "--------", -- 0x372F
        "--------", -- 0x3730
        "--------", -- 0x3731
        "--------", -- 0x3732
        "--------", -- 0x3733
        "--------", -- 0x3734
        "--------", -- 0x3735
        "--------", -- 0x3736
        "--------", -- 0x3737
        "--------", -- 0x3738
        "--------", -- 0x3739
        "--------", -- 0x373A
        "--------", -- 0x373B
        "--------", -- 0x373C
        "--------", -- 0x373D
        "--------", -- 0x373E
        "--------", -- 0x373F
        "--------", -- 0x3740
        "--------", -- 0x3741
        "--------", -- 0x3742
        "--------", -- 0x3743
        "--------", -- 0x3744
        "--------", -- 0x3745
        "--------", -- 0x3746
        "--------", -- 0x3747
        "--------", -- 0x3748
        "--------", -- 0x3749
        "--------", -- 0x374A
        "--------", -- 0x374B
        "--------", -- 0x374C
        "--------", -- 0x374D
        "--------", -- 0x374E
        "--------", -- 0x374F
        "--------", -- 0x3750
        "--------", -- 0x3751
        "--------", -- 0x3752
        "--------", -- 0x3753
        "--------", -- 0x3754
        "--------", -- 0x3755
        "--------", -- 0x3756
        "--------", -- 0x3757
        "--------", -- 0x3758
        "--------", -- 0x3759
        "--------", -- 0x375A
        "--------", -- 0x375B
        "--------", -- 0x375C
        "--------", -- 0x375D
        "--------", -- 0x375E
        "--------", -- 0x375F
        "--------", -- 0x3760
        "--------", -- 0x3761
        "--------", -- 0x3762
        "--------", -- 0x3763
        "--------", -- 0x3764
        "--------", -- 0x3765
        "--------", -- 0x3766
        "--------", -- 0x3767
        "--------", -- 0x3768
        "--------", -- 0x3769
        "--------", -- 0x376A
        "--------", -- 0x376B
        "--------", -- 0x376C
        "--------", -- 0x376D
        "--------", -- 0x376E
        "--------", -- 0x376F
        "--------", -- 0x3770
        "--------", -- 0x3771
        "--------", -- 0x3772
        "--------", -- 0x3773
        "--------", -- 0x3774
        "--------", -- 0x3775
        "--------", -- 0x3776
        "--------", -- 0x3777
        "--------", -- 0x3778
        "--------", -- 0x3779
        "--------", -- 0x377A
        "--------", -- 0x377B
        "--------", -- 0x377C
        "--------", -- 0x377D
        "--------", -- 0x377E
        "--------", -- 0x377F
        "--------", -- 0x3780
        "--------", -- 0x3781
        "--------", -- 0x3782
        "--------", -- 0x3783
        "--------", -- 0x3784
        "--------", -- 0x3785
        "--------", -- 0x3786
        "--------", -- 0x3787
        "--------", -- 0x3788
        "--------", -- 0x3789
        "--------", -- 0x378A
        "--------", -- 0x378B
        "--------", -- 0x378C
        "--------", -- 0x378D
        "--------", -- 0x378E
        "--------", -- 0x378F
        "--------", -- 0x3790
        "--------", -- 0x3791
        "--------", -- 0x3792
        "--------", -- 0x3793
        "--------", -- 0x3794
        "--------", -- 0x3795
        "--------", -- 0x3796
        "--------", -- 0x3797
        "--------", -- 0x3798
        "--------", -- 0x3799
        "--------", -- 0x379A
        "--------", -- 0x379B
        "--------", -- 0x379C
        "--------", -- 0x379D
        "--------", -- 0x379E
        "--------", -- 0x379F
        "--------", -- 0x37A0
        "--------", -- 0x37A1
        "--------", -- 0x37A2
        "--------", -- 0x37A3
        "--------", -- 0x37A4
        "--------", -- 0x37A5
        "--------", -- 0x37A6
        "--------", -- 0x37A7
        "--------", -- 0x37A8
        "--------", -- 0x37A9
        "--------", -- 0x37AA
        "--------", -- 0x37AB
        "--------", -- 0x37AC
        "--------", -- 0x37AD
        "--------", -- 0x37AE
        "--------", -- 0x37AF
        "--------", -- 0x37B0
        "--------", -- 0x37B1
        "--------", -- 0x37B2
        "--------", -- 0x37B3
        "--------", -- 0x37B4
        "--------", -- 0x37B5
        "--------", -- 0x37B6
        "--------", -- 0x37B7
        "--------", -- 0x37B8
        "--------", -- 0x37B9
        "--------", -- 0x37BA
        "--------", -- 0x37BB
        "--------", -- 0x37BC
        "--------", -- 0x37BD
        "--------", -- 0x37BE
        "--------", -- 0x37BF
        "--------", -- 0x37C0
        "--------", -- 0x37C1
        "--------", -- 0x37C2
        "--------", -- 0x37C3
        "--------", -- 0x37C4
        "--------", -- 0x37C5
        "--------", -- 0x37C6
        "--------", -- 0x37C7
        "--------", -- 0x37C8
        "--------", -- 0x37C9
        "--------", -- 0x37CA
        "--------", -- 0x37CB
        "--------", -- 0x37CC
        "--------", -- 0x37CD
        "--------", -- 0x37CE
        "--------", -- 0x37CF
        "--------", -- 0x37D0
        "--------", -- 0x37D1
        "--------", -- 0x37D2
        "--------", -- 0x37D3
        "--------", -- 0x37D4
        "--------", -- 0x37D5
        "--------", -- 0x37D6
        "--------", -- 0x37D7
        "--------", -- 0x37D8
        "--------", -- 0x37D9
        "--------", -- 0x37DA
        "--------", -- 0x37DB
        "--------", -- 0x37DC
        "--------", -- 0x37DD
        "--------", -- 0x37DE
        "--------", -- 0x37DF
        "--------", -- 0x37E0
        "--------", -- 0x37E1
        "--------", -- 0x37E2
        "--------", -- 0x37E3
        "--------", -- 0x37E4
        "--------", -- 0x37E5
        "--------", -- 0x37E6
        "--------", -- 0x37E7
        "--------", -- 0x37E8
        "--------", -- 0x37E9
        "--------", -- 0x37EA
        "--------", -- 0x37EB
        "--------", -- 0x37EC
        "--------", -- 0x37ED
        "--------", -- 0x37EE
        "--------", -- 0x37EF
        "--------", -- 0x37F0
        "--------", -- 0x37F1
        "--------", -- 0x37F2
        "--------", -- 0x37F3
        "--------", -- 0x37F4
        "--------", -- 0x37F5
        "--------", -- 0x37F6
        "--------", -- 0x37F7
        "--------", -- 0x37F8
        "--------", -- 0x37F9
        "--------", -- 0x37FA
        "--------", -- 0x37FB
        "--------", -- 0x37FC
        "--------", -- 0x37FD
        "--------", -- 0x37FE
        "--------", -- 0x37FF
        "--------", -- 0x3800
        "--------", -- 0x3801
        "--------", -- 0x3802
        "--------", -- 0x3803
        "--------", -- 0x3804
        "--------", -- 0x3805
        "--------", -- 0x3806
        "--------", -- 0x3807
        "--------", -- 0x3808
        "--------", -- 0x3809
        "--------", -- 0x380A
        "--------", -- 0x380B
        "--------", -- 0x380C
        "--------", -- 0x380D
        "--------", -- 0x380E
        "--------", -- 0x380F
        "--------", -- 0x3810
        "--------", -- 0x3811
        "--------", -- 0x3812
        "--------", -- 0x3813
        "--------", -- 0x3814
        "--------", -- 0x3815
        "--------", -- 0x3816
        "--------", -- 0x3817
        "--------", -- 0x3818
        "--------", -- 0x3819
        "--------", -- 0x381A
        "--------", -- 0x381B
        "--------", -- 0x381C
        "--------", -- 0x381D
        "--------", -- 0x381E
        "--------", -- 0x381F
        "--------", -- 0x3820
        "--------", -- 0x3821
        "--------", -- 0x3822
        "--------", -- 0x3823
        "--------", -- 0x3824
        "--------", -- 0x3825
        "--------", -- 0x3826
        "--------", -- 0x3827
        "--------", -- 0x3828
        "--------", -- 0x3829
        "--------", -- 0x382A
        "--------", -- 0x382B
        "--------", -- 0x382C
        "--------", -- 0x382D
        "--------", -- 0x382E
        "--------", -- 0x382F
        "--------", -- 0x3830
        "--------", -- 0x3831
        "--------", -- 0x3832
        "--------", -- 0x3833
        "--------", -- 0x3834
        "--------", -- 0x3835
        "--------", -- 0x3836
        "--------", -- 0x3837
        "--------", -- 0x3838
        "--------", -- 0x3839
        "--------", -- 0x383A
        "--------", -- 0x383B
        "--------", -- 0x383C
        "--------", -- 0x383D
        "--------", -- 0x383E
        "--------", -- 0x383F
        "--------", -- 0x3840
        "--------", -- 0x3841
        "--------", -- 0x3842
        "--------", -- 0x3843
        "--------", -- 0x3844
        "--------", -- 0x3845
        "--------", -- 0x3846
        "--------", -- 0x3847
        "--------", -- 0x3848
        "--------", -- 0x3849
        "--------", -- 0x384A
        "--------", -- 0x384B
        "--------", -- 0x384C
        "--------", -- 0x384D
        "--------", -- 0x384E
        "--------", -- 0x384F
        "--------", -- 0x3850
        "--------", -- 0x3851
        "--------", -- 0x3852
        "--------", -- 0x3853
        "--------", -- 0x3854
        "--------", -- 0x3855
        "--------", -- 0x3856
        "--------", -- 0x3857
        "--------", -- 0x3858
        "--------", -- 0x3859
        "--------", -- 0x385A
        "--------", -- 0x385B
        "--------", -- 0x385C
        "--------", -- 0x385D
        "--------", -- 0x385E
        "--------", -- 0x385F
        "--------", -- 0x3860
        "--------", -- 0x3861
        "--------", -- 0x3862
        "--------", -- 0x3863
        "--------", -- 0x3864
        "--------", -- 0x3865
        "--------", -- 0x3866
        "--------", -- 0x3867
        "--------", -- 0x3868
        "--------", -- 0x3869
        "--------", -- 0x386A
        "--------", -- 0x386B
        "--------", -- 0x386C
        "--------", -- 0x386D
        "--------", -- 0x386E
        "--------", -- 0x386F
        "--------", -- 0x3870
        "--------", -- 0x3871
        "--------", -- 0x3872
        "--------", -- 0x3873
        "--------", -- 0x3874
        "--------", -- 0x3875
        "--------", -- 0x3876
        "--------", -- 0x3877
        "--------", -- 0x3878
        "--------", -- 0x3879
        "--------", -- 0x387A
        "--------", -- 0x387B
        "--------", -- 0x387C
        "--------", -- 0x387D
        "--------", -- 0x387E
        "--------", -- 0x387F
        "--------", -- 0x3880
        "--------", -- 0x3881
        "--------", -- 0x3882
        "--------", -- 0x3883
        "--------", -- 0x3884
        "--------", -- 0x3885
        "--------", -- 0x3886
        "--------", -- 0x3887
        "--------", -- 0x3888
        "--------", -- 0x3889
        "--------", -- 0x388A
        "--------", -- 0x388B
        "--------", -- 0x388C
        "--------", -- 0x388D
        "--------", -- 0x388E
        "--------", -- 0x388F
        "--------", -- 0x3890
        "--------", -- 0x3891
        "--------", -- 0x3892
        "--------", -- 0x3893
        "--------", -- 0x3894
        "--------", -- 0x3895
        "--------", -- 0x3896
        "--------", -- 0x3897
        "--------", -- 0x3898
        "--------", -- 0x3899
        "--------", -- 0x389A
        "--------", -- 0x389B
        "--------", -- 0x389C
        "--------", -- 0x389D
        "--------", -- 0x389E
        "--------", -- 0x389F
        "--------", -- 0x38A0
        "--------", -- 0x38A1
        "--------", -- 0x38A2
        "--------", -- 0x38A3
        "--------", -- 0x38A4
        "--------", -- 0x38A5
        "--------", -- 0x38A6
        "--------", -- 0x38A7
        "--------", -- 0x38A8
        "--------", -- 0x38A9
        "--------", -- 0x38AA
        "--------", -- 0x38AB
        "--------", -- 0x38AC
        "--------", -- 0x38AD
        "--------", -- 0x38AE
        "--------", -- 0x38AF
        "--------", -- 0x38B0
        "--------", -- 0x38B1
        "--------", -- 0x38B2
        "--------", -- 0x38B3
        "--------", -- 0x38B4
        "--------", -- 0x38B5
        "--------", -- 0x38B6
        "--------", -- 0x38B7
        "--------", -- 0x38B8
        "--------", -- 0x38B9
        "--------", -- 0x38BA
        "--------", -- 0x38BB
        "--------", -- 0x38BC
        "--------", -- 0x38BD
        "--------", -- 0x38BE
        "--------", -- 0x38BF
        "--------", -- 0x38C0
        "--------", -- 0x38C1
        "--------", -- 0x38C2
        "--------", -- 0x38C3
        "--------", -- 0x38C4
        "--------", -- 0x38C5
        "--------", -- 0x38C6
        "--------", -- 0x38C7
        "--------", -- 0x38C8
        "--------", -- 0x38C9
        "--------", -- 0x38CA
        "--------", -- 0x38CB
        "--------", -- 0x38CC
        "--------", -- 0x38CD
        "--------", -- 0x38CE
        "--------", -- 0x38CF
        "--------", -- 0x38D0
        "--------", -- 0x38D1
        "--------", -- 0x38D2
        "--------", -- 0x38D3
        "--------", -- 0x38D4
        "--------", -- 0x38D5
        "--------", -- 0x38D6
        "--------", -- 0x38D7
        "--------", -- 0x38D8
        "--------", -- 0x38D9
        "--------", -- 0x38DA
        "--------", -- 0x38DB
        "--------", -- 0x38DC
        "--------", -- 0x38DD
        "--------", -- 0x38DE
        "--------", -- 0x38DF
        "--------", -- 0x38E0
        "--------", -- 0x38E1
        "--------", -- 0x38E2
        "--------", -- 0x38E3
        "--------", -- 0x38E4
        "--------", -- 0x38E5
        "--------", -- 0x38E6
        "--------", -- 0x38E7
        "--------", -- 0x38E8
        "--------", -- 0x38E9
        "--------", -- 0x38EA
        "--------", -- 0x38EB
        "--------", -- 0x38EC
        "--------", -- 0x38ED
        "--------", -- 0x38EE
        "--------", -- 0x38EF
        "--------", -- 0x38F0
        "--------", -- 0x38F1
        "--------", -- 0x38F2
        "--------", -- 0x38F3
        "--------", -- 0x38F4
        "--------", -- 0x38F5
        "--------", -- 0x38F6
        "--------", -- 0x38F7
        "--------", -- 0x38F8
        "--------", -- 0x38F9
        "--------", -- 0x38FA
        "--------", -- 0x38FB
        "--------", -- 0x38FC
        "--------", -- 0x38FD
        "--------", -- 0x38FE
        "--------", -- 0x38FF
        "--------", -- 0x3900
        "--------", -- 0x3901
        "--------", -- 0x3902
        "--------", -- 0x3903
        "--------", -- 0x3904
        "--------", -- 0x3905
        "--------", -- 0x3906
        "--------", -- 0x3907
        "--------", -- 0x3908
        "--------", -- 0x3909
        "--------", -- 0x390A
        "--------", -- 0x390B
        "--------", -- 0x390C
        "--------", -- 0x390D
        "--------", -- 0x390E
        "--------", -- 0x390F
        "--------", -- 0x3910
        "--------", -- 0x3911
        "--------", -- 0x3912
        "--------", -- 0x3913
        "--------", -- 0x3914
        "--------", -- 0x3915
        "--------", -- 0x3916
        "--------", -- 0x3917
        "--------", -- 0x3918
        "--------", -- 0x3919
        "--------", -- 0x391A
        "--------", -- 0x391B
        "--------", -- 0x391C
        "--------", -- 0x391D
        "--------", -- 0x391E
        "--------", -- 0x391F
        "--------", -- 0x3920
        "--------", -- 0x3921
        "--------", -- 0x3922
        "--------", -- 0x3923
        "--------", -- 0x3924
        "--------", -- 0x3925
        "--------", -- 0x3926
        "--------", -- 0x3927
        "--------", -- 0x3928
        "--------", -- 0x3929
        "--------", -- 0x392A
        "--------", -- 0x392B
        "--------", -- 0x392C
        "--------", -- 0x392D
        "--------", -- 0x392E
        "--------", -- 0x392F
        "--------", -- 0x3930
        "--------", -- 0x3931
        "--------", -- 0x3932
        "--------", -- 0x3933
        "--------", -- 0x3934
        "--------", -- 0x3935
        "--------", -- 0x3936
        "--------", -- 0x3937
        "--------", -- 0x3938
        "--------", -- 0x3939
        "--------", -- 0x393A
        "--------", -- 0x393B
        "--------", -- 0x393C
        "--------", -- 0x393D
        "--------", -- 0x393E
        "--------", -- 0x393F
        "--------", -- 0x3940
        "--------", -- 0x3941
        "--------", -- 0x3942
        "--------", -- 0x3943
        "--------", -- 0x3944
        "--------", -- 0x3945
        "--------", -- 0x3946
        "--------", -- 0x3947
        "--------", -- 0x3948
        "--------", -- 0x3949
        "--------", -- 0x394A
        "--------", -- 0x394B
        "--------", -- 0x394C
        "--------", -- 0x394D
        "--------", -- 0x394E
        "--------", -- 0x394F
        "--------", -- 0x3950
        "--------", -- 0x3951
        "--------", -- 0x3952
        "--------", -- 0x3953
        "--------", -- 0x3954
        "--------", -- 0x3955
        "--------", -- 0x3956
        "--------", -- 0x3957
        "--------", -- 0x3958
        "--------", -- 0x3959
        "--------", -- 0x395A
        "--------", -- 0x395B
        "--------", -- 0x395C
        "--------", -- 0x395D
        "--------", -- 0x395E
        "--------", -- 0x395F
        "--------", -- 0x3960
        "--------", -- 0x3961
        "--------", -- 0x3962
        "--------", -- 0x3963
        "--------", -- 0x3964
        "--------", -- 0x3965
        "--------", -- 0x3966
        "--------", -- 0x3967
        "--------", -- 0x3968
        "--------", -- 0x3969
        "--------", -- 0x396A
        "--------", -- 0x396B
        "--------", -- 0x396C
        "--------", -- 0x396D
        "--------", -- 0x396E
        "--------", -- 0x396F
        "--------", -- 0x3970
        "--------", -- 0x3971
        "--------", -- 0x3972
        "--------", -- 0x3973
        "--------", -- 0x3974
        "--------", -- 0x3975
        "--------", -- 0x3976
        "--------", -- 0x3977
        "--------", -- 0x3978
        "--------", -- 0x3979
        "--------", -- 0x397A
        "--------", -- 0x397B
        "--------", -- 0x397C
        "--------", -- 0x397D
        "--------", -- 0x397E
        "--------", -- 0x397F
        "--------", -- 0x3980
        "--------", -- 0x3981
        "--------", -- 0x3982
        "--------", -- 0x3983
        "--------", -- 0x3984
        "--------", -- 0x3985
        "--------", -- 0x3986
        "--------", -- 0x3987
        "--------", -- 0x3988
        "--------", -- 0x3989
        "--------", -- 0x398A
        "--------", -- 0x398B
        "--------", -- 0x398C
        "--------", -- 0x398D
        "--------", -- 0x398E
        "--------", -- 0x398F
        "--------", -- 0x3990
        "--------", -- 0x3991
        "--------", -- 0x3992
        "--------", -- 0x3993
        "--------", -- 0x3994
        "--------", -- 0x3995
        "--------", -- 0x3996
        "--------", -- 0x3997
        "--------", -- 0x3998
        "--------", -- 0x3999
        "--------", -- 0x399A
        "--------", -- 0x399B
        "--------", -- 0x399C
        "--------", -- 0x399D
        "--------", -- 0x399E
        "--------", -- 0x399F
        "--------", -- 0x39A0
        "--------", -- 0x39A1
        "--------", -- 0x39A2
        "--------", -- 0x39A3
        "--------", -- 0x39A4
        "--------", -- 0x39A5
        "--------", -- 0x39A6
        "--------", -- 0x39A7
        "--------", -- 0x39A8
        "--------", -- 0x39A9
        "--------", -- 0x39AA
        "--------", -- 0x39AB
        "--------", -- 0x39AC
        "--------", -- 0x39AD
        "--------", -- 0x39AE
        "--------", -- 0x39AF
        "--------", -- 0x39B0
        "--------", -- 0x39B1
        "--------", -- 0x39B2
        "--------", -- 0x39B3
        "--------", -- 0x39B4
        "--------", -- 0x39B5
        "--------", -- 0x39B6
        "--------", -- 0x39B7
        "--------", -- 0x39B8
        "--------", -- 0x39B9
        "--------", -- 0x39BA
        "--------", -- 0x39BB
        "--------", -- 0x39BC
        "--------", -- 0x39BD
        "--------", -- 0x39BE
        "--------", -- 0x39BF
        "--------", -- 0x39C0
        "--------", -- 0x39C1
        "--------", -- 0x39C2
        "--------", -- 0x39C3
        "--------", -- 0x39C4
        "--------", -- 0x39C5
        "--------", -- 0x39C6
        "--------", -- 0x39C7
        "--------", -- 0x39C8
        "--------", -- 0x39C9
        "--------", -- 0x39CA
        "--------", -- 0x39CB
        "--------", -- 0x39CC
        "--------", -- 0x39CD
        "--------", -- 0x39CE
        "--------", -- 0x39CF
        "--------", -- 0x39D0
        "--------", -- 0x39D1
        "--------", -- 0x39D2
        "--------", -- 0x39D3
        "--------", -- 0x39D4
        "--------", -- 0x39D5
        "--------", -- 0x39D6
        "--------", -- 0x39D7
        "--------", -- 0x39D8
        "--------", -- 0x39D9
        "--------", -- 0x39DA
        "--------", -- 0x39DB
        "--------", -- 0x39DC
        "--------", -- 0x39DD
        "--------", -- 0x39DE
        "--------", -- 0x39DF
        "--------", -- 0x39E0
        "--------", -- 0x39E1
        "--------", -- 0x39E2
        "--------", -- 0x39E3
        "--------", -- 0x39E4
        "--------", -- 0x39E5
        "--------", -- 0x39E6
        "--------", -- 0x39E7
        "--------", -- 0x39E8
        "--------", -- 0x39E9
        "--------", -- 0x39EA
        "--------", -- 0x39EB
        "--------", -- 0x39EC
        "--------", -- 0x39ED
        "--------", -- 0x39EE
        "--------", -- 0x39EF
        "--------", -- 0x39F0
        "--------", -- 0x39F1
        "--------", -- 0x39F2
        "--------", -- 0x39F3
        "--------", -- 0x39F4
        "--------", -- 0x39F5
        "--------", -- 0x39F6
        "--------", -- 0x39F7
        "--------", -- 0x39F8
        "--------", -- 0x39F9
        "--------", -- 0x39FA
        "--------", -- 0x39FB
        "--------", -- 0x39FC
        "--------", -- 0x39FD
        "--------", -- 0x39FE
        "--------", -- 0x39FF
        "--------", -- 0x3A00
        "--------", -- 0x3A01
        "--------", -- 0x3A02
        "--------", -- 0x3A03
        "--------", -- 0x3A04
        "--------", -- 0x3A05
        "--------", -- 0x3A06
        "--------", -- 0x3A07
        "--------", -- 0x3A08
        "--------", -- 0x3A09
        "--------", -- 0x3A0A
        "--------", -- 0x3A0B
        "--------", -- 0x3A0C
        "--------", -- 0x3A0D
        "--------", -- 0x3A0E
        "--------", -- 0x3A0F
        "--------", -- 0x3A10
        "--------", -- 0x3A11
        "--------", -- 0x3A12
        "--------", -- 0x3A13
        "--------", -- 0x3A14
        "--------", -- 0x3A15
        "--------", -- 0x3A16
        "--------", -- 0x3A17
        "--------", -- 0x3A18
        "--------", -- 0x3A19
        "--------", -- 0x3A1A
        "--------", -- 0x3A1B
        "--------", -- 0x3A1C
        "--------", -- 0x3A1D
        "--------", -- 0x3A1E
        "--------", -- 0x3A1F
        "--------", -- 0x3A20
        "--------", -- 0x3A21
        "--------", -- 0x3A22
        "--------", -- 0x3A23
        "--------", -- 0x3A24
        "--------", -- 0x3A25
        "--------", -- 0x3A26
        "--------", -- 0x3A27
        "--------", -- 0x3A28
        "--------", -- 0x3A29
        "--------", -- 0x3A2A
        "--------", -- 0x3A2B
        "--------", -- 0x3A2C
        "--------", -- 0x3A2D
        "--------", -- 0x3A2E
        "--------", -- 0x3A2F
        "--------", -- 0x3A30
        "--------", -- 0x3A31
        "--------", -- 0x3A32
        "--------", -- 0x3A33
        "--------", -- 0x3A34
        "--------", -- 0x3A35
        "--------", -- 0x3A36
        "--------", -- 0x3A37
        "--------", -- 0x3A38
        "--------", -- 0x3A39
        "--------", -- 0x3A3A
        "--------", -- 0x3A3B
        "--------", -- 0x3A3C
        "--------", -- 0x3A3D
        "--------", -- 0x3A3E
        "--------", -- 0x3A3F
        "--------", -- 0x3A40
        "--------", -- 0x3A41
        "--------", -- 0x3A42
        "--------", -- 0x3A43
        "--------", -- 0x3A44
        "--------", -- 0x3A45
        "--------", -- 0x3A46
        "--------", -- 0x3A47
        "--------", -- 0x3A48
        "--------", -- 0x3A49
        "--------", -- 0x3A4A
        "--------", -- 0x3A4B
        "--------", -- 0x3A4C
        "--------", -- 0x3A4D
        "--------", -- 0x3A4E
        "--------", -- 0x3A4F
        "--------", -- 0x3A50
        "--------", -- 0x3A51
        "--------", -- 0x3A52
        "--------", -- 0x3A53
        "--------", -- 0x3A54
        "--------", -- 0x3A55
        "--------", -- 0x3A56
        "--------", -- 0x3A57
        "--------", -- 0x3A58
        "--------", -- 0x3A59
        "--------", -- 0x3A5A
        "--------", -- 0x3A5B
        "--------", -- 0x3A5C
        "--------", -- 0x3A5D
        "--------", -- 0x3A5E
        "--------", -- 0x3A5F
        "--------", -- 0x3A60
        "--------", -- 0x3A61
        "--------", -- 0x3A62
        "--------", -- 0x3A63
        "--------", -- 0x3A64
        "--------", -- 0x3A65
        "--------", -- 0x3A66
        "--------", -- 0x3A67
        "--------", -- 0x3A68
        "--------", -- 0x3A69
        "--------", -- 0x3A6A
        "--------", -- 0x3A6B
        "--------", -- 0x3A6C
        "--------", -- 0x3A6D
        "--------", -- 0x3A6E
        "--------", -- 0x3A6F
        "--------", -- 0x3A70
        "--------", -- 0x3A71
        "--------", -- 0x3A72
        "--------", -- 0x3A73
        "--------", -- 0x3A74
        "--------", -- 0x3A75
        "--------", -- 0x3A76
        "--------", -- 0x3A77
        "--------", -- 0x3A78
        "--------", -- 0x3A79
        "--------", -- 0x3A7A
        "--------", -- 0x3A7B
        "--------", -- 0x3A7C
        "--------", -- 0x3A7D
        "--------", -- 0x3A7E
        "--------", -- 0x3A7F
        "--------", -- 0x3A80
        "--------", -- 0x3A81
        "--------", -- 0x3A82
        "--------", -- 0x3A83
        "--------", -- 0x3A84
        "--------", -- 0x3A85
        "--------", -- 0x3A86
        "--------", -- 0x3A87
        "--------", -- 0x3A88
        "--------", -- 0x3A89
        "--------", -- 0x3A8A
        "--------", -- 0x3A8B
        "--------", -- 0x3A8C
        "--------", -- 0x3A8D
        "--------", -- 0x3A8E
        "--------", -- 0x3A8F
        "--------", -- 0x3A90
        "--------", -- 0x3A91
        "--------", -- 0x3A92
        "--------", -- 0x3A93
        "--------", -- 0x3A94
        "--------", -- 0x3A95
        "--------", -- 0x3A96
        "--------", -- 0x3A97
        "--------", -- 0x3A98
        "--------", -- 0x3A99
        "--------", -- 0x3A9A
        "--------", -- 0x3A9B
        "--------", -- 0x3A9C
        "--------", -- 0x3A9D
        "--------", -- 0x3A9E
        "--------", -- 0x3A9F
        "--------", -- 0x3AA0
        "--------", -- 0x3AA1
        "--------", -- 0x3AA2
        "--------", -- 0x3AA3
        "--------", -- 0x3AA4
        "--------", -- 0x3AA5
        "--------", -- 0x3AA6
        "--------", -- 0x3AA7
        "--------", -- 0x3AA8
        "--------", -- 0x3AA9
        "--------", -- 0x3AAA
        "--------", -- 0x3AAB
        "--------", -- 0x3AAC
        "--------", -- 0x3AAD
        "--------", -- 0x3AAE
        "--------", -- 0x3AAF
        "--------", -- 0x3AB0
        "--------", -- 0x3AB1
        "--------", -- 0x3AB2
        "--------", -- 0x3AB3
        "--------", -- 0x3AB4
        "--------", -- 0x3AB5
        "--------", -- 0x3AB6
        "--------", -- 0x3AB7
        "--------", -- 0x3AB8
        "--------", -- 0x3AB9
        "--------", -- 0x3ABA
        "--------", -- 0x3ABB
        "--------", -- 0x3ABC
        "--------", -- 0x3ABD
        "--------", -- 0x3ABE
        "--------", -- 0x3ABF
        "--------", -- 0x3AC0
        "--------", -- 0x3AC1
        "--------", -- 0x3AC2
        "--------", -- 0x3AC3
        "--------", -- 0x3AC4
        "--------", -- 0x3AC5
        "--------", -- 0x3AC6
        "--------", -- 0x3AC7
        "--------", -- 0x3AC8
        "--------", -- 0x3AC9
        "--------", -- 0x3ACA
        "--------", -- 0x3ACB
        "--------", -- 0x3ACC
        "--------", -- 0x3ACD
        "--------", -- 0x3ACE
        "--------", -- 0x3ACF
        "--------", -- 0x3AD0
        "--------", -- 0x3AD1
        "--------", -- 0x3AD2
        "--------", -- 0x3AD3
        "--------", -- 0x3AD4
        "--------", -- 0x3AD5
        "--------", -- 0x3AD6
        "--------", -- 0x3AD7
        "--------", -- 0x3AD8
        "--------", -- 0x3AD9
        "--------", -- 0x3ADA
        "--------", -- 0x3ADB
        "--------", -- 0x3ADC
        "--------", -- 0x3ADD
        "--------", -- 0x3ADE
        "--------", -- 0x3ADF
        "--------", -- 0x3AE0
        "--------", -- 0x3AE1
        "--------", -- 0x3AE2
        "--------", -- 0x3AE3
        "--------", -- 0x3AE4
        "--------", -- 0x3AE5
        "--------", -- 0x3AE6
        "--------", -- 0x3AE7
        "--------", -- 0x3AE8
        "--------", -- 0x3AE9
        "--------", -- 0x3AEA
        "--------", -- 0x3AEB
        "--------", -- 0x3AEC
        "--------", -- 0x3AED
        "--------", -- 0x3AEE
        "--------", -- 0x3AEF
        "--------", -- 0x3AF0
        "--------", -- 0x3AF1
        "--------", -- 0x3AF2
        "--------", -- 0x3AF3
        "--------", -- 0x3AF4
        "--------", -- 0x3AF5
        "--------", -- 0x3AF6
        "--------", -- 0x3AF7
        "--------", -- 0x3AF8
        "--------", -- 0x3AF9
        "--------", -- 0x3AFA
        "--------", -- 0x3AFB
        "--------", -- 0x3AFC
        "--------", -- 0x3AFD
        "--------", -- 0x3AFE
        "--------", -- 0x3AFF
        "--------", -- 0x3B00
        "--------", -- 0x3B01
        "--------", -- 0x3B02
        "--------", -- 0x3B03
        "--------", -- 0x3B04
        "--------", -- 0x3B05
        "--------", -- 0x3B06
        "--------", -- 0x3B07
        "--------", -- 0x3B08
        "--------", -- 0x3B09
        "--------", -- 0x3B0A
        "--------", -- 0x3B0B
        "--------", -- 0x3B0C
        "--------", -- 0x3B0D
        "--------", -- 0x3B0E
        "--------", -- 0x3B0F
        "--------", -- 0x3B10
        "--------", -- 0x3B11
        "--------", -- 0x3B12
        "--------", -- 0x3B13
        "--------", -- 0x3B14
        "--------", -- 0x3B15
        "--------", -- 0x3B16
        "--------", -- 0x3B17
        "--------", -- 0x3B18
        "--------", -- 0x3B19
        "--------", -- 0x3B1A
        "--------", -- 0x3B1B
        "--------", -- 0x3B1C
        "--------", -- 0x3B1D
        "--------", -- 0x3B1E
        "--------", -- 0x3B1F
        "--------", -- 0x3B20
        "--------", -- 0x3B21
        "--------", -- 0x3B22
        "--------", -- 0x3B23
        "--------", -- 0x3B24
        "--------", -- 0x3B25
        "--------", -- 0x3B26
        "--------", -- 0x3B27
        "--------", -- 0x3B28
        "--------", -- 0x3B29
        "--------", -- 0x3B2A
        "--------", -- 0x3B2B
        "--------", -- 0x3B2C
        "--------", -- 0x3B2D
        "--------", -- 0x3B2E
        "--------", -- 0x3B2F
        "--------", -- 0x3B30
        "--------", -- 0x3B31
        "--------", -- 0x3B32
        "--------", -- 0x3B33
        "--------", -- 0x3B34
        "--------", -- 0x3B35
        "--------", -- 0x3B36
        "--------", -- 0x3B37
        "--------", -- 0x3B38
        "--------", -- 0x3B39
        "--------", -- 0x3B3A
        "--------", -- 0x3B3B
        "--------", -- 0x3B3C
        "--------", -- 0x3B3D
        "--------", -- 0x3B3E
        "--------", -- 0x3B3F
        "--------", -- 0x3B40
        "--------", -- 0x3B41
        "--------", -- 0x3B42
        "--------", -- 0x3B43
        "--------", -- 0x3B44
        "--------", -- 0x3B45
        "--------", -- 0x3B46
        "--------", -- 0x3B47
        "--------", -- 0x3B48
        "--------", -- 0x3B49
        "--------", -- 0x3B4A
        "--------", -- 0x3B4B
        "--------", -- 0x3B4C
        "--------", -- 0x3B4D
        "--------", -- 0x3B4E
        "--------", -- 0x3B4F
        "--------", -- 0x3B50
        "--------", -- 0x3B51
        "--------", -- 0x3B52
        "--------", -- 0x3B53
        "--------", -- 0x3B54
        "--------", -- 0x3B55
        "--------", -- 0x3B56
        "--------", -- 0x3B57
        "--------", -- 0x3B58
        "--------", -- 0x3B59
        "--------", -- 0x3B5A
        "--------", -- 0x3B5B
        "--------", -- 0x3B5C
        "--------", -- 0x3B5D
        "--------", -- 0x3B5E
        "--------", -- 0x3B5F
        "--------", -- 0x3B60
        "--------", -- 0x3B61
        "--------", -- 0x3B62
        "--------", -- 0x3B63
        "--------", -- 0x3B64
        "--------", -- 0x3B65
        "--------", -- 0x3B66
        "--------", -- 0x3B67
        "--------", -- 0x3B68
        "--------", -- 0x3B69
        "--------", -- 0x3B6A
        "--------", -- 0x3B6B
        "--------", -- 0x3B6C
        "--------", -- 0x3B6D
        "--------", -- 0x3B6E
        "--------", -- 0x3B6F
        "--------", -- 0x3B70
        "--------", -- 0x3B71
        "--------", -- 0x3B72
        "--------", -- 0x3B73
        "--------", -- 0x3B74
        "--------", -- 0x3B75
        "--------", -- 0x3B76
        "--------", -- 0x3B77
        "--------", -- 0x3B78
        "--------", -- 0x3B79
        "--------", -- 0x3B7A
        "--------", -- 0x3B7B
        "--------", -- 0x3B7C
        "--------", -- 0x3B7D
        "--------", -- 0x3B7E
        "--------", -- 0x3B7F
        "--------", -- 0x3B80
        "--------", -- 0x3B81
        "--------", -- 0x3B82
        "--------", -- 0x3B83
        "--------", -- 0x3B84
        "--------", -- 0x3B85
        "--------", -- 0x3B86
        "--------", -- 0x3B87
        "--------", -- 0x3B88
        "--------", -- 0x3B89
        "--------", -- 0x3B8A
        "--------", -- 0x3B8B
        "--------", -- 0x3B8C
        "--------", -- 0x3B8D
        "--------", -- 0x3B8E
        "--------", -- 0x3B8F
        "--------", -- 0x3B90
        "--------", -- 0x3B91
        "--------", -- 0x3B92
        "--------", -- 0x3B93
        "--------", -- 0x3B94
        "--------", -- 0x3B95
        "--------", -- 0x3B96
        "--------", -- 0x3B97
        "--------", -- 0x3B98
        "--------", -- 0x3B99
        "--------", -- 0x3B9A
        "--------", -- 0x3B9B
        "--------", -- 0x3B9C
        "--------", -- 0x3B9D
        "--------", -- 0x3B9E
        "--------", -- 0x3B9F
        "--------", -- 0x3BA0
        "--------", -- 0x3BA1
        "--------", -- 0x3BA2
        "--------", -- 0x3BA3
        "--------", -- 0x3BA4
        "--------", -- 0x3BA5
        "--------", -- 0x3BA6
        "--------", -- 0x3BA7
        "--------", -- 0x3BA8
        "--------", -- 0x3BA9
        "--------", -- 0x3BAA
        "--------", -- 0x3BAB
        "--------", -- 0x3BAC
        "--------", -- 0x3BAD
        "--------", -- 0x3BAE
        "--------", -- 0x3BAF
        "--------", -- 0x3BB0
        "--------", -- 0x3BB1
        "--------", -- 0x3BB2
        "--------", -- 0x3BB3
        "--------", -- 0x3BB4
        "--------", -- 0x3BB5
        "--------", -- 0x3BB6
        "--------", -- 0x3BB7
        "--------", -- 0x3BB8
        "--------", -- 0x3BB9
        "--------", -- 0x3BBA
        "--------", -- 0x3BBB
        "--------", -- 0x3BBC
        "--------", -- 0x3BBD
        "--------", -- 0x3BBE
        "--------", -- 0x3BBF
        "--------", -- 0x3BC0
        "--------", -- 0x3BC1
        "--------", -- 0x3BC2
        "--------", -- 0x3BC3
        "--------", -- 0x3BC4
        "--------", -- 0x3BC5
        "--------", -- 0x3BC6
        "--------", -- 0x3BC7
        "--------", -- 0x3BC8
        "--------", -- 0x3BC9
        "--------", -- 0x3BCA
        "--------", -- 0x3BCB
        "--------", -- 0x3BCC
        "--------", -- 0x3BCD
        "--------", -- 0x3BCE
        "--------", -- 0x3BCF
        "--------", -- 0x3BD0
        "--------", -- 0x3BD1
        "--------", -- 0x3BD2
        "--------", -- 0x3BD3
        "--------", -- 0x3BD4
        "--------", -- 0x3BD5
        "--------", -- 0x3BD6
        "--------", -- 0x3BD7
        "--------", -- 0x3BD8
        "--------", -- 0x3BD9
        "--------", -- 0x3BDA
        "--------", -- 0x3BDB
        "--------", -- 0x3BDC
        "--------", -- 0x3BDD
        "--------", -- 0x3BDE
        "--------", -- 0x3BDF
        "--------", -- 0x3BE0
        "--------", -- 0x3BE1
        "--------", -- 0x3BE2
        "--------", -- 0x3BE3
        "--------", -- 0x3BE4
        "--------", -- 0x3BE5
        "--------", -- 0x3BE6
        "--------", -- 0x3BE7
        "--------", -- 0x3BE8
        "--------", -- 0x3BE9
        "--------", -- 0x3BEA
        "--------", -- 0x3BEB
        "--------", -- 0x3BEC
        "--------", -- 0x3BED
        "--------", -- 0x3BEE
        "--------", -- 0x3BEF
        "--------", -- 0x3BF0
        "--------", -- 0x3BF1
        "--------", -- 0x3BF2
        "--------", -- 0x3BF3
        "--------", -- 0x3BF4
        "--------", -- 0x3BF5
        "--------", -- 0x3BF6
        "--------", -- 0x3BF7
        "--------", -- 0x3BF8
        "--------", -- 0x3BF9
        "--------", -- 0x3BFA
        "--------", -- 0x3BFB
        "--------", -- 0x3BFC
        "--------", -- 0x3BFD
        "--------", -- 0x3BFE
        "--------", -- 0x3BFF
        "--------", -- 0x3C00
        "--------", -- 0x3C01
        "--------", -- 0x3C02
        "--------", -- 0x3C03
        "--------", -- 0x3C04
        "--------", -- 0x3C05
        "--------", -- 0x3C06
        "--------", -- 0x3C07
        "--------", -- 0x3C08
        "--------", -- 0x3C09
        "--------", -- 0x3C0A
        "--------", -- 0x3C0B
        "--------", -- 0x3C0C
        "--------", -- 0x3C0D
        "--------", -- 0x3C0E
        "--------", -- 0x3C0F
        "--------", -- 0x3C10
        "--------", -- 0x3C11
        "--------", -- 0x3C12
        "--------", -- 0x3C13
        "--------", -- 0x3C14
        "--------", -- 0x3C15
        "--------", -- 0x3C16
        "--------", -- 0x3C17
        "--------", -- 0x3C18
        "--------", -- 0x3C19
        "--------", -- 0x3C1A
        "--------", -- 0x3C1B
        "--------", -- 0x3C1C
        "--------", -- 0x3C1D
        "--------", -- 0x3C1E
        "--------", -- 0x3C1F
        "--------", -- 0x3C20
        "--------", -- 0x3C21
        "--------", -- 0x3C22
        "--------", -- 0x3C23
        "--------", -- 0x3C24
        "--------", -- 0x3C25
        "--------", -- 0x3C26
        "--------", -- 0x3C27
        "--------", -- 0x3C28
        "--------", -- 0x3C29
        "--------", -- 0x3C2A
        "--------", -- 0x3C2B
        "--------", -- 0x3C2C
        "--------", -- 0x3C2D
        "--------", -- 0x3C2E
        "--------", -- 0x3C2F
        "--------", -- 0x3C30
        "--------", -- 0x3C31
        "--------", -- 0x3C32
        "--------", -- 0x3C33
        "--------", -- 0x3C34
        "--------", -- 0x3C35
        "--------", -- 0x3C36
        "--------", -- 0x3C37
        "--------", -- 0x3C38
        "--------", -- 0x3C39
        "--------", -- 0x3C3A
        "--------", -- 0x3C3B
        "--------", -- 0x3C3C
        "--------", -- 0x3C3D
        "--------", -- 0x3C3E
        "--------", -- 0x3C3F
        "--------", -- 0x3C40
        "--------", -- 0x3C41
        "--------", -- 0x3C42
        "--------", -- 0x3C43
        "--------", -- 0x3C44
        "--------", -- 0x3C45
        "--------", -- 0x3C46
        "--------", -- 0x3C47
        "--------", -- 0x3C48
        "--------", -- 0x3C49
        "--------", -- 0x3C4A
        "--------", -- 0x3C4B
        "--------", -- 0x3C4C
        "--------", -- 0x3C4D
        "--------", -- 0x3C4E
        "--------", -- 0x3C4F
        "--------", -- 0x3C50
        "--------", -- 0x3C51
        "--------", -- 0x3C52
        "--------", -- 0x3C53
        "--------", -- 0x3C54
        "--------", -- 0x3C55
        "--------", -- 0x3C56
        "--------", -- 0x3C57
        "--------", -- 0x3C58
        "--------", -- 0x3C59
        "--------", -- 0x3C5A
        "--------", -- 0x3C5B
        "--------", -- 0x3C5C
        "--------", -- 0x3C5D
        "--------", -- 0x3C5E
        "--------", -- 0x3C5F
        "--------", -- 0x3C60
        "--------", -- 0x3C61
        "--------", -- 0x3C62
        "--------", -- 0x3C63
        "--------", -- 0x3C64
        "--------", -- 0x3C65
        "--------", -- 0x3C66
        "--------", -- 0x3C67
        "--------", -- 0x3C68
        "--------", -- 0x3C69
        "--------", -- 0x3C6A
        "--------", -- 0x3C6B
        "--------", -- 0x3C6C
        "--------", -- 0x3C6D
        "--------", -- 0x3C6E
        "--------", -- 0x3C6F
        "--------", -- 0x3C70
        "--------", -- 0x3C71
        "--------", -- 0x3C72
        "--------", -- 0x3C73
        "--------", -- 0x3C74
        "--------", -- 0x3C75
        "--------", -- 0x3C76
        "--------", -- 0x3C77
        "--------", -- 0x3C78
        "--------", -- 0x3C79
        "--------", -- 0x3C7A
        "--------", -- 0x3C7B
        "--------", -- 0x3C7C
        "--------", -- 0x3C7D
        "--------", -- 0x3C7E
        "--------", -- 0x3C7F
        "--------", -- 0x3C80
        "--------", -- 0x3C81
        "--------", -- 0x3C82
        "--------", -- 0x3C83
        "--------", -- 0x3C84
        "--------", -- 0x3C85
        "--------", -- 0x3C86
        "--------", -- 0x3C87
        "--------", -- 0x3C88
        "--------", -- 0x3C89
        "--------", -- 0x3C8A
        "--------", -- 0x3C8B
        "--------", -- 0x3C8C
        "--------", -- 0x3C8D
        "--------", -- 0x3C8E
        "--------", -- 0x3C8F
        "--------", -- 0x3C90
        "--------", -- 0x3C91
        "--------", -- 0x3C92
        "--------", -- 0x3C93
        "--------", -- 0x3C94
        "--------", -- 0x3C95
        "--------", -- 0x3C96
        "--------", -- 0x3C97
        "--------", -- 0x3C98
        "--------", -- 0x3C99
        "--------", -- 0x3C9A
        "--------", -- 0x3C9B
        "--------", -- 0x3C9C
        "--------", -- 0x3C9D
        "--------", -- 0x3C9E
        "--------", -- 0x3C9F
        "--------", -- 0x3CA0
        "--------", -- 0x3CA1
        "--------", -- 0x3CA2
        "--------", -- 0x3CA3
        "--------", -- 0x3CA4
        "--------", -- 0x3CA5
        "--------", -- 0x3CA6
        "--------", -- 0x3CA7
        "--------", -- 0x3CA8
        "--------", -- 0x3CA9
        "--------", -- 0x3CAA
        "--------", -- 0x3CAB
        "--------", -- 0x3CAC
        "--------", -- 0x3CAD
        "--------", -- 0x3CAE
        "--------", -- 0x3CAF
        "--------", -- 0x3CB0
        "--------", -- 0x3CB1
        "--------", -- 0x3CB2
        "--------", -- 0x3CB3
        "--------", -- 0x3CB4
        "--------", -- 0x3CB5
        "--------", -- 0x3CB6
        "--------", -- 0x3CB7
        "--------", -- 0x3CB8
        "--------", -- 0x3CB9
        "--------", -- 0x3CBA
        "--------", -- 0x3CBB
        "--------", -- 0x3CBC
        "--------", -- 0x3CBD
        "--------", -- 0x3CBE
        "--------", -- 0x3CBF
        "--------", -- 0x3CC0
        "--------", -- 0x3CC1
        "--------", -- 0x3CC2
        "--------", -- 0x3CC3
        "--------", -- 0x3CC4
        "--------", -- 0x3CC5
        "--------", -- 0x3CC6
        "--------", -- 0x3CC7
        "--------", -- 0x3CC8
        "--------", -- 0x3CC9
        "--------", -- 0x3CCA
        "--------", -- 0x3CCB
        "--------", -- 0x3CCC
        "--------", -- 0x3CCD
        "--------", -- 0x3CCE
        "--------", -- 0x3CCF
        "--------", -- 0x3CD0
        "--------", -- 0x3CD1
        "--------", -- 0x3CD2
        "--------", -- 0x3CD3
        "--------", -- 0x3CD4
        "--------", -- 0x3CD5
        "--------", -- 0x3CD6
        "--------", -- 0x3CD7
        "--------", -- 0x3CD8
        "--------", -- 0x3CD9
        "--------", -- 0x3CDA
        "--------", -- 0x3CDB
        "--------", -- 0x3CDC
        "--------", -- 0x3CDD
        "--------", -- 0x3CDE
        "--------", -- 0x3CDF
        "--------", -- 0x3CE0
        "--------", -- 0x3CE1
        "--------", -- 0x3CE2
        "--------", -- 0x3CE3
        "--------", -- 0x3CE4
        "--------", -- 0x3CE5
        "--------", -- 0x3CE6
        "--------", -- 0x3CE7
        "--------", -- 0x3CE8
        "--------", -- 0x3CE9
        "--------", -- 0x3CEA
        "--------", -- 0x3CEB
        "--------", -- 0x3CEC
        "--------", -- 0x3CED
        "--------", -- 0x3CEE
        "--------", -- 0x3CEF
        "--------", -- 0x3CF0
        "--------", -- 0x3CF1
        "--------", -- 0x3CF2
        "--------", -- 0x3CF3
        "--------", -- 0x3CF4
        "--------", -- 0x3CF5
        "--------", -- 0x3CF6
        "--------", -- 0x3CF7
        "--------", -- 0x3CF8
        "--------", -- 0x3CF9
        "--------", -- 0x3CFA
        "--------", -- 0x3CFB
        "--------", -- 0x3CFC
        "--------", -- 0x3CFD
        "--------", -- 0x3CFE
        "--------", -- 0x3CFF
        "--------", -- 0x3D00
        "--------", -- 0x3D01
        "--------", -- 0x3D02
        "--------", -- 0x3D03
        "--------", -- 0x3D04
        "--------", -- 0x3D05
        "--------", -- 0x3D06
        "--------", -- 0x3D07
        "--------", -- 0x3D08
        "--------", -- 0x3D09
        "--------", -- 0x3D0A
        "--------", -- 0x3D0B
        "--------", -- 0x3D0C
        "--------", -- 0x3D0D
        "--------", -- 0x3D0E
        "--------", -- 0x3D0F
        "--------", -- 0x3D10
        "--------", -- 0x3D11
        "--------", -- 0x3D12
        "--------", -- 0x3D13
        "--------", -- 0x3D14
        "--------", -- 0x3D15
        "--------", -- 0x3D16
        "--------", -- 0x3D17
        "--------", -- 0x3D18
        "--------", -- 0x3D19
        "--------", -- 0x3D1A
        "--------", -- 0x3D1B
        "--------", -- 0x3D1C
        "--------", -- 0x3D1D
        "--------", -- 0x3D1E
        "--------", -- 0x3D1F
        "--------", -- 0x3D20
        "--------", -- 0x3D21
        "--------", -- 0x3D22
        "--------", -- 0x3D23
        "--------", -- 0x3D24
        "--------", -- 0x3D25
        "--------", -- 0x3D26
        "--------", -- 0x3D27
        "--------", -- 0x3D28
        "--------", -- 0x3D29
        "--------", -- 0x3D2A
        "--------", -- 0x3D2B
        "--------", -- 0x3D2C
        "--------", -- 0x3D2D
        "--------", -- 0x3D2E
        "--------", -- 0x3D2F
        "--------", -- 0x3D30
        "--------", -- 0x3D31
        "--------", -- 0x3D32
        "--------", -- 0x3D33
        "--------", -- 0x3D34
        "--------", -- 0x3D35
        "--------", -- 0x3D36
        "--------", -- 0x3D37
        "--------", -- 0x3D38
        "--------", -- 0x3D39
        "--------", -- 0x3D3A
        "--------", -- 0x3D3B
        "--------", -- 0x3D3C
        "--------", -- 0x3D3D
        "--------", -- 0x3D3E
        "--------", -- 0x3D3F
        "--------", -- 0x3D40
        "--------", -- 0x3D41
        "--------", -- 0x3D42
        "--------", -- 0x3D43
        "--------", -- 0x3D44
        "--------", -- 0x3D45
        "--------", -- 0x3D46
        "--------", -- 0x3D47
        "--------", -- 0x3D48
        "--------", -- 0x3D49
        "--------", -- 0x3D4A
        "--------", -- 0x3D4B
        "--------", -- 0x3D4C
        "--------", -- 0x3D4D
        "--------", -- 0x3D4E
        "--------", -- 0x3D4F
        "--------", -- 0x3D50
        "--------", -- 0x3D51
        "--------", -- 0x3D52
        "--------", -- 0x3D53
        "--------", -- 0x3D54
        "--------", -- 0x3D55
        "--------", -- 0x3D56
        "--------", -- 0x3D57
        "--------", -- 0x3D58
        "--------", -- 0x3D59
        "--------", -- 0x3D5A
        "--------", -- 0x3D5B
        "--------", -- 0x3D5C
        "--------", -- 0x3D5D
        "--------", -- 0x3D5E
        "--------", -- 0x3D5F
        "--------", -- 0x3D60
        "--------", -- 0x3D61
        "--------", -- 0x3D62
        "--------", -- 0x3D63
        "--------", -- 0x3D64
        "--------", -- 0x3D65
        "--------", -- 0x3D66
        "--------", -- 0x3D67
        "--------", -- 0x3D68
        "--------", -- 0x3D69
        "--------", -- 0x3D6A
        "--------", -- 0x3D6B
        "--------", -- 0x3D6C
        "--------", -- 0x3D6D
        "--------", -- 0x3D6E
        "--------", -- 0x3D6F
        "--------", -- 0x3D70
        "--------", -- 0x3D71
        "--------", -- 0x3D72
        "--------", -- 0x3D73
        "--------", -- 0x3D74
        "--------", -- 0x3D75
        "--------", -- 0x3D76
        "--------", -- 0x3D77
        "--------", -- 0x3D78
        "--------", -- 0x3D79
        "--------", -- 0x3D7A
        "--------", -- 0x3D7B
        "--------", -- 0x3D7C
        "--------", -- 0x3D7D
        "--------", -- 0x3D7E
        "--------", -- 0x3D7F
        "--------", -- 0x3D80
        "--------", -- 0x3D81
        "--------", -- 0x3D82
        "--------", -- 0x3D83
        "--------", -- 0x3D84
        "--------", -- 0x3D85
        "--------", -- 0x3D86
        "--------", -- 0x3D87
        "--------", -- 0x3D88
        "--------", -- 0x3D89
        "--------", -- 0x3D8A
        "--------", -- 0x3D8B
        "--------", -- 0x3D8C
        "--------", -- 0x3D8D
        "--------", -- 0x3D8E
        "--------", -- 0x3D8F
        "--------", -- 0x3D90
        "--------", -- 0x3D91
        "--------", -- 0x3D92
        "--------", -- 0x3D93
        "--------", -- 0x3D94
        "--------", -- 0x3D95
        "--------", -- 0x3D96
        "--------", -- 0x3D97
        "--------", -- 0x3D98
        "--------", -- 0x3D99
        "--------", -- 0x3D9A
        "--------", -- 0x3D9B
        "--------", -- 0x3D9C
        "--------", -- 0x3D9D
        "--------", -- 0x3D9E
        "--------", -- 0x3D9F
        "--------", -- 0x3DA0
        "--------", -- 0x3DA1
        "--------", -- 0x3DA2
        "--------", -- 0x3DA3
        "--------", -- 0x3DA4
        "--------", -- 0x3DA5
        "--------", -- 0x3DA6
        "--------", -- 0x3DA7
        "--------", -- 0x3DA8
        "--------", -- 0x3DA9
        "--------", -- 0x3DAA
        "--------", -- 0x3DAB
        "--------", -- 0x3DAC
        "--------", -- 0x3DAD
        "--------", -- 0x3DAE
        "--------", -- 0x3DAF
        "--------", -- 0x3DB0
        "--------", -- 0x3DB1
        "--------", -- 0x3DB2
        "--------", -- 0x3DB3
        "--------", -- 0x3DB4
        "--------", -- 0x3DB5
        "--------", -- 0x3DB6
        "--------", -- 0x3DB7
        "--------", -- 0x3DB8
        "--------", -- 0x3DB9
        "--------", -- 0x3DBA
        "--------", -- 0x3DBB
        "--------", -- 0x3DBC
        "--------", -- 0x3DBD
        "--------", -- 0x3DBE
        "--------", -- 0x3DBF
        "--------", -- 0x3DC0
        "--------", -- 0x3DC1
        "--------", -- 0x3DC2
        "--------", -- 0x3DC3
        "--------", -- 0x3DC4
        "--------", -- 0x3DC5
        "--------", -- 0x3DC6
        "--------", -- 0x3DC7
        "--------", -- 0x3DC8
        "--------", -- 0x3DC9
        "--------", -- 0x3DCA
        "--------", -- 0x3DCB
        "--------", -- 0x3DCC
        "--------", -- 0x3DCD
        "--------", -- 0x3DCE
        "--------", -- 0x3DCF
        "--------", -- 0x3DD0
        "--------", -- 0x3DD1
        "--------", -- 0x3DD2
        "--------", -- 0x3DD3
        "--------", -- 0x3DD4
        "--------", -- 0x3DD5
        "--------", -- 0x3DD6
        "--------", -- 0x3DD7
        "--------", -- 0x3DD8
        "--------", -- 0x3DD9
        "--------", -- 0x3DDA
        "--------", -- 0x3DDB
        "--------", -- 0x3DDC
        "--------", -- 0x3DDD
        "--------", -- 0x3DDE
        "--------", -- 0x3DDF
        "--------", -- 0x3DE0
        "--------", -- 0x3DE1
        "--------", -- 0x3DE2
        "--------", -- 0x3DE3
        "--------", -- 0x3DE4
        "--------", -- 0x3DE5
        "--------", -- 0x3DE6
        "--------", -- 0x3DE7
        "--------", -- 0x3DE8
        "--------", -- 0x3DE9
        "--------", -- 0x3DEA
        "--------", -- 0x3DEB
        "--------", -- 0x3DEC
        "--------", -- 0x3DED
        "--------", -- 0x3DEE
        "--------", -- 0x3DEF
        "--------", -- 0x3DF0
        "--------", -- 0x3DF1
        "--------", -- 0x3DF2
        "--------", -- 0x3DF3
        "--------", -- 0x3DF4
        "--------", -- 0x3DF5
        "--------", -- 0x3DF6
        "--------", -- 0x3DF7
        "--------", -- 0x3DF8
        "--------", -- 0x3DF9
        "--------", -- 0x3DFA
        "--------", -- 0x3DFB
        "--------", -- 0x3DFC
        "--------", -- 0x3DFD
        "--------", -- 0x3DFE
        "--------", -- 0x3DFF
        "--------", -- 0x3E00
        "--------", -- 0x3E01
        "--------", -- 0x3E02
        "--------", -- 0x3E03
        "--------", -- 0x3E04
        "--------", -- 0x3E05
        "--------", -- 0x3E06
        "--------", -- 0x3E07
        "--------", -- 0x3E08
        "--------", -- 0x3E09
        "--------", -- 0x3E0A
        "--------", -- 0x3E0B
        "--------", -- 0x3E0C
        "--------", -- 0x3E0D
        "--------", -- 0x3E0E
        "--------", -- 0x3E0F
        "--------", -- 0x3E10
        "--------", -- 0x3E11
        "--------", -- 0x3E12
        "--------", -- 0x3E13
        "--------", -- 0x3E14
        "--------", -- 0x3E15
        "--------", -- 0x3E16
        "--------", -- 0x3E17
        "--------", -- 0x3E18
        "--------", -- 0x3E19
        "--------", -- 0x3E1A
        "--------", -- 0x3E1B
        "--------", -- 0x3E1C
        "--------", -- 0x3E1D
        "--------", -- 0x3E1E
        "--------", -- 0x3E1F
        "--------", -- 0x3E20
        "--------", -- 0x3E21
        "--------", -- 0x3E22
        "--------", -- 0x3E23
        "--------", -- 0x3E24
        "--------", -- 0x3E25
        "--------", -- 0x3E26
        "--------", -- 0x3E27
        "--------", -- 0x3E28
        "--------", -- 0x3E29
        "--------", -- 0x3E2A
        "--------", -- 0x3E2B
        "--------", -- 0x3E2C
        "--------", -- 0x3E2D
        "--------", -- 0x3E2E
        "--------", -- 0x3E2F
        "--------", -- 0x3E30
        "--------", -- 0x3E31
        "--------", -- 0x3E32
        "--------", -- 0x3E33
        "--------", -- 0x3E34
        "--------", -- 0x3E35
        "--------", -- 0x3E36
        "--------", -- 0x3E37
        "--------", -- 0x3E38
        "--------", -- 0x3E39
        "--------", -- 0x3E3A
        "--------", -- 0x3E3B
        "--------", -- 0x3E3C
        "--------", -- 0x3E3D
        "--------", -- 0x3E3E
        "--------", -- 0x3E3F
        "--------", -- 0x3E40
        "--------", -- 0x3E41
        "--------", -- 0x3E42
        "--------", -- 0x3E43
        "--------", -- 0x3E44
        "--------", -- 0x3E45
        "--------", -- 0x3E46
        "--------", -- 0x3E47
        "--------", -- 0x3E48
        "--------", -- 0x3E49
        "--------", -- 0x3E4A
        "--------", -- 0x3E4B
        "--------", -- 0x3E4C
        "--------", -- 0x3E4D
        "--------", -- 0x3E4E
        "--------", -- 0x3E4F
        "--------", -- 0x3E50
        "--------", -- 0x3E51
        "--------", -- 0x3E52
        "--------", -- 0x3E53
        "--------", -- 0x3E54
        "--------", -- 0x3E55
        "--------", -- 0x3E56
        "--------", -- 0x3E57
        "--------", -- 0x3E58
        "--------", -- 0x3E59
        "--------", -- 0x3E5A
        "--------", -- 0x3E5B
        "--------", -- 0x3E5C
        "--------", -- 0x3E5D
        "--------", -- 0x3E5E
        "--------", -- 0x3E5F
        "--------", -- 0x3E60
        "--------", -- 0x3E61
        "--------", -- 0x3E62
        "--------", -- 0x3E63
        "--------", -- 0x3E64
        "--------", -- 0x3E65
        "--------", -- 0x3E66
        "--------", -- 0x3E67
        "--------", -- 0x3E68
        "--------", -- 0x3E69
        "--------", -- 0x3E6A
        "--------", -- 0x3E6B
        "--------", -- 0x3E6C
        "--------", -- 0x3E6D
        "--------", -- 0x3E6E
        "--------", -- 0x3E6F
        "--------", -- 0x3E70
        "--------", -- 0x3E71
        "--------", -- 0x3E72
        "--------", -- 0x3E73
        "--------", -- 0x3E74
        "--------", -- 0x3E75
        "--------", -- 0x3E76
        "--------", -- 0x3E77
        "--------", -- 0x3E78
        "--------", -- 0x3E79
        "--------", -- 0x3E7A
        "--------", -- 0x3E7B
        "--------", -- 0x3E7C
        "--------", -- 0x3E7D
        "--------", -- 0x3E7E
        "--------", -- 0x3E7F
        "--------", -- 0x3E80
        "--------", -- 0x3E81
        "--------", -- 0x3E82
        "--------", -- 0x3E83
        "--------", -- 0x3E84
        "--------", -- 0x3E85
        "--------", -- 0x3E86
        "--------", -- 0x3E87
        "--------", -- 0x3E88
        "--------", -- 0x3E89
        "--------", -- 0x3E8A
        "--------", -- 0x3E8B
        "--------", -- 0x3E8C
        "--------", -- 0x3E8D
        "--------", -- 0x3E8E
        "--------", -- 0x3E8F
        "--------", -- 0x3E90
        "--------", -- 0x3E91
        "--------", -- 0x3E92
        "--------", -- 0x3E93
        "--------", -- 0x3E94
        "--------", -- 0x3E95
        "--------", -- 0x3E96
        "--------", -- 0x3E97
        "--------", -- 0x3E98
        "--------", -- 0x3E99
        "--------", -- 0x3E9A
        "--------", -- 0x3E9B
        "--------", -- 0x3E9C
        "--------", -- 0x3E9D
        "--------", -- 0x3E9E
        "--------", -- 0x3E9F
        "--------", -- 0x3EA0
        "--------", -- 0x3EA1
        "--------", -- 0x3EA2
        "--------", -- 0x3EA3
        "--------", -- 0x3EA4
        "--------", -- 0x3EA5
        "--------", -- 0x3EA6
        "--------", -- 0x3EA7
        "--------", -- 0x3EA8
        "--------", -- 0x3EA9
        "--------", -- 0x3EAA
        "--------", -- 0x3EAB
        "--------", -- 0x3EAC
        "--------", -- 0x3EAD
        "--------", -- 0x3EAE
        "--------", -- 0x3EAF
        "--------", -- 0x3EB0
        "--------", -- 0x3EB1
        "--------", -- 0x3EB2
        "--------", -- 0x3EB3
        "--------", -- 0x3EB4
        "--------", -- 0x3EB5
        "--------", -- 0x3EB6
        "--------", -- 0x3EB7
        "--------", -- 0x3EB8
        "--------", -- 0x3EB9
        "--------", -- 0x3EBA
        "--------", -- 0x3EBB
        "--------", -- 0x3EBC
        "--------", -- 0x3EBD
        "--------", -- 0x3EBE
        "--------", -- 0x3EBF
        "--------", -- 0x3EC0
        "--------", -- 0x3EC1
        "--------", -- 0x3EC2
        "--------", -- 0x3EC3
        "--------", -- 0x3EC4
        "--------", -- 0x3EC5
        "--------", -- 0x3EC6
        "--------", -- 0x3EC7
        "--------", -- 0x3EC8
        "--------", -- 0x3EC9
        "--------", -- 0x3ECA
        "--------", -- 0x3ECB
        "--------", -- 0x3ECC
        "--------", -- 0x3ECD
        "--------", -- 0x3ECE
        "--------", -- 0x3ECF
        "--------", -- 0x3ED0
        "--------", -- 0x3ED1
        "--------", -- 0x3ED2
        "--------", -- 0x3ED3
        "--------", -- 0x3ED4
        "--------", -- 0x3ED5
        "--------", -- 0x3ED6
        "--------", -- 0x3ED7
        "--------", -- 0x3ED8
        "--------", -- 0x3ED9
        "--------", -- 0x3EDA
        "--------", -- 0x3EDB
        "--------", -- 0x3EDC
        "--------", -- 0x3EDD
        "--------", -- 0x3EDE
        "--------", -- 0x3EDF
        "--------", -- 0x3EE0
        "--------", -- 0x3EE1
        "--------", -- 0x3EE2
        "--------", -- 0x3EE3
        "--------", -- 0x3EE4
        "--------", -- 0x3EE5
        "--------", -- 0x3EE6
        "--------", -- 0x3EE7
        "--------", -- 0x3EE8
        "--------", -- 0x3EE9
        "--------", -- 0x3EEA
        "--------", -- 0x3EEB
        "--------", -- 0x3EEC
        "--------", -- 0x3EED
        "--------", -- 0x3EEE
        "--------", -- 0x3EEF
        "--------", -- 0x3EF0
        "--------", -- 0x3EF1
        "--------", -- 0x3EF2
        "--------", -- 0x3EF3
        "--------", -- 0x3EF4
        "--------", -- 0x3EF5
        "--------", -- 0x3EF6
        "--------", -- 0x3EF7
        "--------", -- 0x3EF8
        "--------", -- 0x3EF9
        "--------", -- 0x3EFA
        "--------", -- 0x3EFB
        "--------", -- 0x3EFC
        "--------", -- 0x3EFD
        "--------", -- 0x3EFE
        "--------", -- 0x3EFF
        "--------", -- 0x3F00
        "--------", -- 0x3F01
        "--------", -- 0x3F02
        "--------", -- 0x3F03
        "--------", -- 0x3F04
        "--------", -- 0x3F05
        "--------", -- 0x3F06
        "--------", -- 0x3F07
        "--------", -- 0x3F08
        "--------", -- 0x3F09
        "--------", -- 0x3F0A
        "--------", -- 0x3F0B
        "--------", -- 0x3F0C
        "--------", -- 0x3F0D
        "--------", -- 0x3F0E
        "--------", -- 0x3F0F
        "--------", -- 0x3F10
        "--------", -- 0x3F11
        "--------", -- 0x3F12
        "--------", -- 0x3F13
        "--------", -- 0x3F14
        "--------", -- 0x3F15
        "--------", -- 0x3F16
        "--------", -- 0x3F17
        "--------", -- 0x3F18
        "--------", -- 0x3F19
        "--------", -- 0x3F1A
        "--------", -- 0x3F1B
        "--------", -- 0x3F1C
        "--------", -- 0x3F1D
        "--------", -- 0x3F1E
        "--------", -- 0x3F1F
        "--------", -- 0x3F20
        "--------", -- 0x3F21
        "--------", -- 0x3F22
        "--------", -- 0x3F23
        "--------", -- 0x3F24
        "--------", -- 0x3F25
        "--------", -- 0x3F26
        "--------", -- 0x3F27
        "--------", -- 0x3F28
        "--------", -- 0x3F29
        "--------", -- 0x3F2A
        "--------", -- 0x3F2B
        "--------", -- 0x3F2C
        "--------", -- 0x3F2D
        "--------", -- 0x3F2E
        "--------", -- 0x3F2F
        "--------", -- 0x3F30
        "--------", -- 0x3F31
        "--------", -- 0x3F32
        "--------", -- 0x3F33
        "--------", -- 0x3F34
        "--------", -- 0x3F35
        "--------", -- 0x3F36
        "--------", -- 0x3F37
        "--------", -- 0x3F38
        "--------", -- 0x3F39
        "--------", -- 0x3F3A
        "--------", -- 0x3F3B
        "--------", -- 0x3F3C
        "--------", -- 0x3F3D
        "--------", -- 0x3F3E
        "--------", -- 0x3F3F
        "--------", -- 0x3F40
        "--------", -- 0x3F41
        "--------", -- 0x3F42
        "--------", -- 0x3F43
        "--------", -- 0x3F44
        "--------", -- 0x3F45
        "--------", -- 0x3F46
        "--------", -- 0x3F47
        "--------", -- 0x3F48
        "--------", -- 0x3F49
        "--------", -- 0x3F4A
        "--------", -- 0x3F4B
        "--------", -- 0x3F4C
        "--------", -- 0x3F4D
        "--------", -- 0x3F4E
        "--------", -- 0x3F4F
        "--------", -- 0x3F50
        "--------", -- 0x3F51
        "--------", -- 0x3F52
        "--------", -- 0x3F53
        "--------", -- 0x3F54
        "--------", -- 0x3F55
        "--------", -- 0x3F56
        "--------", -- 0x3F57
        "--------", -- 0x3F58
        "--------", -- 0x3F59
        "--------", -- 0x3F5A
        "--------", -- 0x3F5B
        "--------", -- 0x3F5C
        "--------", -- 0x3F5D
        "--------", -- 0x3F5E
        "--------", -- 0x3F5F
        "--------", -- 0x3F60
        "--------", -- 0x3F61
        "--------", -- 0x3F62
        "--------", -- 0x3F63
        "--------", -- 0x3F64
        "--------", -- 0x3F65
        "--------", -- 0x3F66
        "--------", -- 0x3F67
        "--------", -- 0x3F68
        "--------", -- 0x3F69
        "--------", -- 0x3F6A
        "--------", -- 0x3F6B
        "--------", -- 0x3F6C
        "--------", -- 0x3F6D
        "--------", -- 0x3F6E
        "--------", -- 0x3F6F
        "--------", -- 0x3F70
        "--------", -- 0x3F71
        "--------", -- 0x3F72
        "--------", -- 0x3F73
        "--------", -- 0x3F74
        "--------", -- 0x3F75
        "--------", -- 0x3F76
        "--------", -- 0x3F77
        "--------", -- 0x3F78
        "--------", -- 0x3F79
        "--------", -- 0x3F7A
        "--------", -- 0x3F7B
        "--------", -- 0x3F7C
        "--------", -- 0x3F7D
        "--------", -- 0x3F7E
        "--------", -- 0x3F7F
        "--------", -- 0x3F80
        "--------", -- 0x3F81
        "--------", -- 0x3F82
        "--------", -- 0x3F83
        "--------", -- 0x3F84
        "--------", -- 0x3F85
        "--------", -- 0x3F86
        "--------", -- 0x3F87
        "--------", -- 0x3F88
        "--------", -- 0x3F89
        "--------", -- 0x3F8A
        "--------", -- 0x3F8B
        "--------", -- 0x3F8C
        "--------", -- 0x3F8D
        "--------", -- 0x3F8E
        "--------", -- 0x3F8F
        "--------", -- 0x3F90
        "--------", -- 0x3F91
        "--------", -- 0x3F92
        "--------", -- 0x3F93
        "--------", -- 0x3F94
        "--------", -- 0x3F95
        "--------", -- 0x3F96
        "--------", -- 0x3F97
        "--------", -- 0x3F98
        "--------", -- 0x3F99
        "--------", -- 0x3F9A
        "--------", -- 0x3F9B
        "--------", -- 0x3F9C
        "--------", -- 0x3F9D
        "--------", -- 0x3F9E
        "--------", -- 0x3F9F
        "--------", -- 0x3FA0
        "--------", -- 0x3FA1
        "--------", -- 0x3FA2
        "--------", -- 0x3FA3
        "--------", -- 0x3FA4
        "--------", -- 0x3FA5
        "--------", -- 0x3FA6
        "--------", -- 0x3FA7
        "--------", -- 0x3FA8
        "--------", -- 0x3FA9
        "--------", -- 0x3FAA
        "--------", -- 0x3FAB
        "--------", -- 0x3FAC
        "--------", -- 0x3FAD
        "--------", -- 0x3FAE
        "--------", -- 0x3FAF
        "--------", -- 0x3FB0
        "--------", -- 0x3FB1
        "--------", -- 0x3FB2
        "--------", -- 0x3FB3
        "--------", -- 0x3FB4
        "--------", -- 0x3FB5
        "--------", -- 0x3FB6
        "--------", -- 0x3FB7
        "--------", -- 0x3FB8
        "--------", -- 0x3FB9
        "--------", -- 0x3FBA
        "--------", -- 0x3FBB
        "--------", -- 0x3FBC
        "--------", -- 0x3FBD
        "--------", -- 0x3FBE
        "--------", -- 0x3FBF
        "--------", -- 0x3FC0
        "--------", -- 0x3FC1
        "--------", -- 0x3FC2
        "--------", -- 0x3FC3
        "--------", -- 0x3FC4
        "--------", -- 0x3FC5
        "--------", -- 0x3FC6
        "--------", -- 0x3FC7
        "--------", -- 0x3FC8
        "--------", -- 0x3FC9
        "--------", -- 0x3FCA
        "--------", -- 0x3FCB
        "--------", -- 0x3FCC
        "--------", -- 0x3FCD
        "--------", -- 0x3FCE
        "--------", -- 0x3FCF
        "--------", -- 0x3FD0
        "--------", -- 0x3FD1
        "--------", -- 0x3FD2
        "--------", -- 0x3FD3
        "--------", -- 0x3FD4
        "--------", -- 0x3FD5
        "--------", -- 0x3FD6
        "--------", -- 0x3FD7
        "--------", -- 0x3FD8
        "--------", -- 0x3FD9
        "--------", -- 0x3FDA
        "--------", -- 0x3FDB
        "--------", -- 0x3FDC
        "--------", -- 0x3FDD
        "--------", -- 0x3FDE
        "--------", -- 0x3FDF
        "--------", -- 0x3FE0
        "--------", -- 0x3FE1
        "--------", -- 0x3FE2
        "--------", -- 0x3FE3
        "--------", -- 0x3FE4
        "--------", -- 0x3FE5
        "--------", -- 0x3FE6
        "--------", -- 0x3FE7
        "--------", -- 0x3FE8
        "--------", -- 0x3FE9
        "--------", -- 0x3FEA
        "--------", -- 0x3FEB
        "--------", -- 0x3FEC
        "--------", -- 0x3FED
        "--------", -- 0x3FEE
        "--------", -- 0x3FEF
        "--------", -- 0x3FF0
        "--------", -- 0x3FF1
        "--------", -- 0x3FF2
        "--------", -- 0x3FF3
        "--------", -- 0x3FF4
        "--------", -- 0x3FF5
        "--------", -- 0x3FF6
        "--------", -- 0x3FF7
        "--------", -- 0x3FF8
        "--------", -- 0x3FF9
        "--------", -- 0x3FFA
        "--------", -- 0x3FFB
        "--------", -- 0x3FFC
        "--------", -- 0x3FFD
        "--------", -- 0x3FFE
        "--------");    -- 0x3FFF
begin
    D <= ROM(to_integer(unsigned(A)));
end;

