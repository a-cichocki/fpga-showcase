--------------------------------------------------------------------------------
-- Project           :  STIX/IDPU/EM
-- Drawing           :  
-- File title        :  
-- Design unit name  :  Stix_pkg
-- Authors           :  A. Cichocki
-- Company           :  Centrum Badañ Kosmicznych
-- Current revision  :  1 (2016-09-27)
--------------------------------------------------------------------------------
-- Description       : 
--------------------------------------------------------------------------------
-- Generated By XmlOutGen v. 1.26
--------------------------------------------------------------------------------

library Cbk;
    use Cbk.DetCtrl_pkg.all;

library grlib;
    use grlib.amba.all;

library ieee;
    use ieee.std_logic_1164.all;

library techmap;
    use techmap.gencomp.all;


package Stix_pkg is 
    type IdefxEvent_t is record
        AsicAddr                                               : std_logic_vector(4 downto 0);
        AdcVal                                                 : std_logic_vector(31 downto 0);
        Strobe                                                 : std_logic;
    end record;
    type IdefxCmdIn_t is record
        CmdStb                                                 : std_logic;
        GrpAddr                                                : std_logic_vector(3 downto 0);
        ReadMode                                               : std_logic_vector(15 downto 0);
        CmdCounter                                             : std_logic_vector(3 downto 0);
        Enable                                                 : std_logic_vector(15 downto 0);
        CmdData                                                : std_logic_vector(15 downto 0);
        WriteMask                                              : std_logic_vector(15 downto 0);
        DelayModeAdc                                           : std_logic_vector(1 downto 0);
        TLatency                                               : std_logic_vector(3 downto 0);
        DelayModeIdefx                                         : std_logic_vector(1 downto 0);
    end record;
    type IdefxCmdOut_t is record
        CmdReady                                               : std_logic;
        ResponseData                                           : std_logic_vector(15 downto 0);
        CmdCounter                                             : std_logic_vector(3 downto 0);
        CmdData                                                : std_logic_vector(15 downto 0);
        GrpAddr                                                : std_logic_vector(3 downto 0);
    end record;
    type ReadoutFsmIn_t is record
        Reset                                                  : std_logic;
        IntegrationTimeMin                                     : std_logic_vector(15 downto 0);
        CalDmask                                               : std_logic_vector(31 downto 0);
        IntegrationTimeMax                                     : std_logic_vector(15 downto 0);
        IntegrationEventsMax                                   : std_logic_vector(31 downto 0);
        ActiveTlut                                             : std_logic;
        CalTq                                                  : std_logic_vector(15 downto 0);
        QlIntTime                                              : std_logic_vector(15 downto 0);
        SetCalEnable                                           : std_logic;
        CalClear                                               : std_logic;
        Wstb                                                   : std_logic;
        SetEnable                                              : std_logic;
        ClearEnable                                            : std_logic;
        QlClear                                                : std_logic;
        CalIrqEn                                               : std_logic;
        QlIrqEn                                                : std_logic;
        FifoIrqEn                                              : std_logic;
        OverflowClear                                          : std_logic;
        QlVarEMask                                             : std_logic_vector(31 downto 0);
        QlVarDMask                                             : std_logic_vector(31 downto 0);
        QlVarPMask                                             : std_logic_vector(11 downto 0);
        SumDMask                                               : std_logic_vector(31 downto 0);
        SumEMask                                               : std_logic_vector(31 downto 0);
    end record;
    type ReadoutFsmOut_t is record
        GroupAddr                                              : std_logic_vector(3 downto 0);
        PixelAddr                                              : std_logic_vector(3 downto 0);
        AsicAddr                                               : std_logic;
        AdcVal                                                 : std_logic_vector(11 downto 0);
        AdcCorVal                                              : std_logic_vector(11 downto 0);
        Energy                                                 : std_logic_vector(4 downto 0);
        Overflow                                               : std_logic;
        EventCount                                             : std_logic_vector(31 downto 0);
        Irq                                                    : std_logic;
        ActiveQL                                               : std_logic_vector(1 downto 0);
        ActiveNominal                                          : std_logic;
        CalCount                                               : std_logic_vector(31 downto 0);
        CalTruncate                                            : std_logic_vector(20 downto 0);
        QlReady                                                : std_logic;
        Enable                                                 : std_logic;
        CalReady                                               : std_logic;
        CalEnable                                              : std_logic;
    end record;
    type QuarterCtrlIn_t is record
        Power                                                  : std_logic_vector(3 downto 0);
        TestPulse                                              : std_logic;
        DacVal                                                 : std_logic_vector(11 downto 0);
        PulseMask                                              : std_logic_vector(3 downto 0);
    end record;
    type QuarterCtrlOut_t is record
        Seu                                                    : std_logic_vector(3 downto 0);
        PulseBusy                                              : std_logic;
        DacVal                                                 : std_logic_vector(11 downto 0);
        PulseMask                                              : std_logic_vector(3 downto 0);
    end record;
    type QuarterIn_t is record
        POWERON                                                : std_logic;
        DACDIN                                                 : std_logic;
        DACSCLK                                                : std_logic;
        DACSYNC_N                                              : std_logic;
        TESTPULSE                                              : std_logic;
    end record;
    type QuarterOut_t is record
        Seu                                                    : std_logic;
    end record;
    type DetGrpIn_t is record
        DinEn                                                  : std_logic;
        Din                                                    : std_logic;
        Stb                                                    : std_logic;
        AdcSclk                                                : std_logic;
        AdcCs                                                  : std_logic;
    end record;
    type DetGrpOut_t is record
        Dout                                                   : std_logic;
        AdcDout                                                : std_logic;
    end record;
    type RotbDetIn_t is record
        ActiveNominal                                          : std_logic;
        ActiveQl                                               : std_logic_vector(1 downto 0);
    end record;
    type ApbRotbOut_t is record
        TestMode                                               : std_logic;
        EdacOn                                                 : std_logic;
        RefreshRate                                            : std_logic_vector(7 downto 0);
        ScrubRate                                              : std_logic_vector(1 downto 0);
        Command                                                : std_logic_vector(1 downto 0);
        EdacReset                                              : std_logic;
        CmdStrobe                                              : std_logic;
        Enable                                                 : std_logic;
    end record;
    type ApbRotbIn_t is record
        SecCount                                               : std_logic_vector(7 downto 0);
        Ready                                                  : std_logic;
        DeDetected                                             : std_logic;
        BlockCount                                             : std_logic_vector(16 downto 0);
        Full                                                   : std_logic;
        Irq                                                    : std_logic;
        IrqSd                                                  : std_logic;
    end record;
    type RotbAsOut_t is record
        Rd                                                     : std_logic;
        Addr                                                   : std_logic_vector(7 downto 0);
    end record;
    type RotbAsIn_t is record
        Data                                                   : std_logic_vector(15 downto 0);
        DataPartition                                          : std_logic;
    end record;
    type CacheRotbIn_t is record
        Address                                                : std_logic_vector(20 downto 0);
        Rd                                                     : std_logic;
    end record;
    type CacheRotbOut_t is record
        Data                                                   : std_logic_vector(31 downto 0);
        Ready                                                  : std_logic;
    end record;
    type AhbRotbIn_t is record
        Ready                                                  : std_logic;
        Data                                                   : std_logic_vector(31 downto 0);
    end record;
    type AhbRotbOut_t is record
        Address                                                : std_logic_vector(6 downto 0);
        Data                                                   : std_logic_vector(31 downto 0);
        Wr                                                     : std_logic;
        Rd                                                     : std_logic;
    end record;
    subtype HkThreshold_t is std_logic_vector(11 downto 0);
    type AspHkIn_t is record
        READ                                                   : std_logic;
        TEMPADDR                                               : std_logic_vector(3 downto 0);
    end record;
    type AspHkOut_t is record
        READY                                                  : std_logic_vector(1 downto 0);
        VAL                                                    : std_logic_vector(11 downto 0);
    end record;
    type ApbAsOut_t is record
        AOn                                                    : std_logic;
        BOn                                                    : std_logic;
        AvgSize                                                : std_logic_vector(2 downto 0);
    end record;
    subtype AspDiodeData_t is std_logic_vector(15 downto 0);
    type ApbTimerIn_t is record
        SubSecond                                              : std_logic_vector(15 downto 0);
        Seconds                                                : std_logic_vector(31 downto 0);
    end record;
    type ApbTimerOut_t is record
        SubSecond                                              : std_logic_vector(15 downto 0);
        Seconds                                                : std_logic_vector(31 downto 0);
        SubSecWstb                                             : std_logic;
    end record;
    type ApbAttnOut_t is record
        SlowRampTimeQuant                                      : std_logic_vector(11 downto 0);
        FastRampTimeQuant                                      : std_logic_vector(7 downto 0);
        Command                                                : std_logic_vector(3 downto 0);
        CmdStrobe                                              : std_logic;
        PWMConfigStrobe1                                       : std_logic;
        ErrorMask                                              : std_logic;
    end record;
    type ApbAttnIn_t is record
        PositionAb                                             : std_logic;
        PositionBc                                             : std_logic;
        Timeout                                                : std_logic;
        Motor1Used                                             : std_logic;
        Motor2Used                                             : std_logic;
        OperationStatus                                        : std_logic;
        SlowRampTimeQuant                                      : std_logic_vector(11 downto 0);
        FastRampTimeQuant                                      : std_logic_vector(7 downto 0);
        ErrorMask                                              : std_logic;
        FailFlag                                               : std_logic;
    end record;
    type CacheDetOut_t is record
        SramDout                                               : std_logic_vector(31 downto 0);
        Bram1Dout                                              : std_logic_vector(15 downto 0);
        Bram4Dout                                              : std_logic_vector(23 downto 0);
        BramTrigDout                                           : std_logic_vector(23 downto 0);
        SramReady                                              : std_logic;
        Bram1Ready                                             : std_logic;
        Bram4Ready                                             : std_logic;
        BramTrigReady                                          : std_logic;
    end record;
    type CacheDetIn_t is record
        SramDin                                                : std_logic_vector(31 downto 0);
        SramAddr                                               : std_logic_vector(18 downto 0);
        SramWr                                                 : std_logic;
        SramRd                                                 : std_logic;
        Bram1Din                                               : std_logic_vector(15 downto 0);
        Bram1Addr                                              : std_logic_vector(7 downto 0);
        Bram1Wr                                                : std_logic;
        Bram1Rd                                                : std_logic;
        Bram4Din                                               : std_logic_vector(23 downto 0);
        Bram4Addr                                              : std_logic_vector(5 downto 0);
        Bram4Wr                                                : std_logic;
        Bram4Rd                                                : std_logic;
        BramTrigDin                                            : std_logic_vector(23 downto 0);
        BramTrigAddr                                           : std_logic_vector(4 downto 0);
        BramTrigWr                                             : std_logic;
        BramTrigRd                                             : std_logic;
    end record;
    type ApbCacheOut_t is record
        OpMode                                                 : std_logic;
        ScrubRate                                              : std_logic_vector(1 downto 0);
        EdacOn                                                 : std_logic;
        EdacReset                                              : std_logic;
        Strobe                                                 : std_logic;
    end record;
    type ApbCacheIn_t is record
        SecCount                                               : std_logic_vector(7 downto 0);
        DeDetected                                             : std_logic;
        Irq                                                    : std_logic;
    end record;
    type AhbCacheOut_t is record
        Address                                                : std_logic_vector(20 downto 0);
        Data                                                   : std_logic_vector(31 downto 0);
        Wr                                                     : std_logic;
        Rd                                                     : std_logic;
    end record;
    type AhbCacheIn_t is record
        Ready                                                  : std_logic;
        Data                                                   : std_logic_vector(31 downto 0);
        Ded                                                    : std_logic;
    end record;
    type ApbGenRegOut_t is record
        WriteStrobe                                            : std_logic;
        CleanShutDown                                          : std_logic;
        StatusClear                                            : std_logic;
        RotbEnabled                                            : std_logic;
        Magic                                                  : std_logic_vector(31 downto 0);
        MagicWStb                                              : std_logic;
        WdogWstb                                               : std_logic;
        WdogCmd                                                : std_logic_vector(2 downto 0);
        WdogReload                                             : std_logic_vector(5 downto 0);
        TickEnabled                                            : std_logic;
    end record;
    type ApbGenRegIn_t is record
        CleanShutDown                                          : std_logic;
        HwRelease                                              : std_logic_vector(5 downto 0);
        HwBuild                                                : std_logic_vector(15 downto 0);
        ThisIdpu                                               : std_logic;
        OtherIsOn                                              : std_logic;
        WatchDog                                               : std_logic;
        Irq                                                    : std_logic;
        Magic                                                  : std_logic_vector(31 downto 0);
        WdogCount                                              : std_logic_vector(5 downto 0);
        WdogReload                                             : std_logic_vector(5 downto 0);
    end record;
    type IdefxEventVector_t is array (15 downto 0) of IdefxEvent_t;
    type ApbDetOut_t is record
        ReadoutFsm                                             : ReadoutFsmIn_t;
        QuarterCtrl                                            : QuarterCtrlIn_t;
        IdefxCtrls                                             : IdefxCmdIn_t;
        SeuIrqEn                                               : std_logic_vector(3 downto 0);
    end record;
    type ApbDetIn_t is record
        ReadoutFsm                                             : ReadoutFsmOut_t;
        QuarterCtrl                                            : QuarterCtrlOut_t;
        IdefxResponse                                          : IdefxCmdOut_t;
        Irq                                                    : std_logic;
    end record;
    type QuarterInVector_t is array (1 to 4) of QuarterIn_t;
    type QuarterOutVector_t is array (1 to 4) of QuarterOut_t;
    type DetGrpInVector_t is array (1 to 16) of DetGrpIn_t;
    type DetGrpOutVector_t is array (1 to 16) of DetGrpOut_t;
    type HkThresholdVector_t is array (1 to 9) of HkThreshold_t;
    type AspQlData_t is array (1 to 4) of AspDiodeData_t;
    type DetPinOut_t is record
        Quarters                                               : QuarterInVector_t;
        DetGrps                                                : DetGrpInVector_t;
    end record;
    type DetPinIn_t is record
        Quarters                                               : QuarterOutVector_t;
        DetGrps                                                : DetGrpOutVector_t;
    end record;
    type ApbHkOut_t is record
        LvEn                                                   : std_logic;
        Hv0116en                                               : std_logic;
        Hv1732en                                               : std_logic;
        AdcAddress                                             : std_logic_vector(6 downto 0);
        Hv0116val                                              : std_logic_vector(7 downto 0);
        Hv1732val                                              : std_logic_vector(7 downto 0);
        Thresholds                                             : HkThresholdVector_t;
        Token                                                  : std_logic_vector(7 downto 0);
        ProtEn                                                 : std_logic_vector(1 to 9);
        IrqEn                                                  : std_logic_vector(1 to 9);
        SpwEn                                                  : std_logic_vector(1 downto 0);
        ThreshWrStb                                            : std_logic_vector(1 to 9);
        TokenWrStb                                             : std_logic;
        ProtClear                                              : std_logic_vector(1 to 9);
    end record;
    type ApbHkIn_t is record
        ProtStat                                               : std_logic_vector(1 to 9);
        AdcReady                                               : std_logic;
        AdcVal                                                 : std_logic_vector(11 downto 0);
        Irq                                                    : std_logic;
        PowerStat                                              : std_logic_vector(4 downto 0);
        ProtEn                                                 : std_logic_vector(1 to 9);
        Thresholds                                             : HkThresholdVector_t;
        BadSample                                              : std_logic_vector(11 downto 0);
    end record;
    type ApbAsIn_t is record
        QlData                                                 : AspQlData_t;
    end record;
    component AdcConfig is 
        port (
            iClk                                                   : in std_logic;
            iRst_n                                                 : in std_logic;
            iAdcEn                                                 : in std_logic;
            iDout                                                  : in std_logic;
            oSclk                                                  : out std_logic;
            oIrq                                                   : out std_logic;
            oData                                                  : out std_logic_vector(15 downto 0);
            iTick                                                  : in std_logic
        );
    end component;
    component IdefxConfig is 
        generic (
            Technology                                             : integer;
            ADC_CS_N_POL                                           : std_logic
        );
        port (
            iClk                                                   : in std_logic;
            iRst_n                                                 : in std_logic;
            iIdefxDout                                             : in std_logic;
            oIdefxDin                                              : out std_logic;
            oIdefxStb                                              : out std_logic;
            iCmdStb                                                : in std_logic;
            iCmdData                                               : in std_logic_vector(15 downto 0);
            iCmdCounter                                            : in std_logic_vector(3 downto 0);
            oReadData                                              : out std_logic_vector(15 downto 0);
            oCmdRdy                                                : out std_logic;
            oAdcSclk                                               : out std_logic;
            oAdcCs_n                                               : out std_logic;
            iAdcDout                                               : in std_logic
        );
    end component;
    component IdefxClkGen is 
        generic (
            ADC_CS_N_POL                                           : std_logic;
            STB_LEN_BITS                                           : integer;
            T_LEN_BITS                                             : integer;
            STB_LEN                                                : integer;
            T_BUFF_LEN                                             : integer;
            T_MUX_LEN                                              : integer;
            T_SETTLE_LEN                                           : integer;
            T_RESET_LEN                                            : integer;
            Technology                                             : integer
        );
        port (
            iClk                                                   : in std_logic;
            iRst_N                                                 : in std_logic;
            oIdefxStb                                              : out std_logic;
            oAdcCs_n                                               : out std_logic;
            oAdcSclkMask                                           : out std_logic;
            oAdcGo                                                 : out std_logic;
            iTLatency                                              : in std_logic_vector(3 downto 0);
            iAdcIrq                                                : in std_logic;
            oIdefxDinEn                                            : out std_logic;
            iEnable                                                : in std_logic;
            iIdefxDout                                             : in std_logic;
            oBusy                                                  : out std_logic;
            iDelayMode                                             : in std_logic_vector(1 downto 0);
            oIrq                                                   : out std_logic;
            oIdefxAddr                                             : out std_logic_vector(4 downto 0);
            oIdefxDin                                              : out std_logic
        );
    end component;
    component AdcIdefxRead is 
        generic (
            ADC_SCLK_LEN_BITS                                      : integer;
            ADC_SCLK_LEN                                           : integer
        );
        port (
            iClk                                                   : in std_logic;
            iRst_N                                                 : in std_logic;
            iAdcGo                                                 : in std_logic;
            oAdcSclk                                               : out std_logic;
            iAdcDout                                               : in std_logic;
            oAdcData                                               : out std_logic_vector(31 downto 0);
            oAdcIrq                                                : out std_logic;
            iDelayMode                                             : in std_logic_vector(1 downto 0)
        );
    end component;
    component Idefx is 
        generic (
            Technology                                             : integer;
            ADC_CS_N_POL                                           : std_logic;
            STB_LEN_BITS                                           : integer;
            T_LEN_BITS                                             : integer;
            STB_LEN                                                : integer;
            T_BUFF_LEN                                             : integer;
            T_MUX_LEN                                              : integer;
            T_SETTLE_LEN                                           : integer;
            T_RESET_LEN                                            : integer;
            ADC_SCLK_LEN_BITS                                      : integer;
            ADC_SCLK_LEN                                           : integer
        );
        port (
            iClk                                                   : in std_logic;
            iRst_n                                                 : in std_logic;
            iEnable                                                : in std_logic;
            iTLatency                                              : in std_logic_vector(3 downto 0);
            oIdefxStb                                              : out std_logic;
            oIdefxDin                                              : out std_logic;
            oIdefxDinEn                                            : out std_logic;
            iIdefxDout                                             : in std_logic;
            oAdcCs                                                 : out std_logic;
            oAdcSclk                                               : out std_logic;
            iAdcDout                                               : in std_logic;
            oIdefxAddr                                             : out std_logic_vector(4 downto 0);
            oAdcData                                               : out std_logic_vector(31 downto 0);
            oIrq                                                   : out std_logic;
            oBusy                                                  : out std_logic;
            iDelayModeAdc                                          : in std_logic_vector(1 downto 0);
            iDelayModeIdefx                                        : in std_logic_vector(1 downto 0)
        );
    end component;
    component IdefxCtrls is 
        generic (
            Technology                                             : integer;
            ADC_CS_N_POL                                           : std_logic;
            STB_LEN_BITS                                           : integer;
            T_LEN_BITS                                             : integer;
            STB_LEN                                                : integer;
            T_BUFF_LEN                                             : integer;
            T_MUX_LEN                                              : integer;
            T_SETTLE_LEN                                           : integer;
            T_RESET_LEN                                            : integer;
            ADC_SCLK_LEN_BITS                                      : integer;
            ADC_SCLK_LEN                                           : integer
        );
        port (
            oEvents                                                : out IdefxEventVector_t;
            iCmd                                                   : in IdefxCmdIn_t;
            oCmd                                                   : out IdefxCmdOut_t;
            iClkF                                                  : in std_logic;
            iRstF_n                                                : in std_logic;
            iDetGrps                                               : in DetGrpOutVector_t;
            oDetGrps                                               : out DetGrpInVector_t;
            iClkM                                                  : in std_logic;
            iRstM_n                                                : in std_logic
        );
    end component;
    component FifoLogic is 
        generic (
            N                                                      : integer;
            Technology                                             : integer
        );
        port (
            iClk                                                   : in std_logic;
            iRst_n                                                 : in std_logic;
            iPush                                                  : in std_logic;
            iPop                                                   : in std_logic;
            iInit                                                  : in std_logic;
            oAdd_w                                                 : out std_logic_vector(N-1 downto 0);
            oAdd_r                                                 : out std_logic_vector(N-1 downto 0);
            oFull                                                  : out std_logic;
            oEmpty                                                 : out std_logic;
            oWe                                                    : out std_logic;
            oRe                                                    : out std_logic;
            oOverFlow                                              : out std_logic;
            oNoPop                                                 : out std_logic
        );
    end component;
    component Fifo is 
        generic (
            Technology                                             : integer;
            N                                                      : integer;
            W                                                      : integer
        );
        port (
            iClk                                                   : in std_logic;
            iRst_n                                                 : in std_logic;
            iPush                                                  : in std_logic;
            iPop                                                   : in std_logic;
            iInit                                                  : in std_logic;
            iDin                                                   : in std_logic_vector(W-1 downto 0);
            oDout                                                  : out std_logic_vector(W-1 downto 0);
            oFull                                                  : out std_logic;
            oEmpty                                                 : out std_logic;
            oOverFlow                                              : out std_logic;
            oNoPop                                                 : out std_logic
        );
    end component;
    component EventReader is 
        port (
            iClk                                                   : in std_logic;
            iRst_n                                                 : in std_logic;
            iEnable                                                : in std_logic;
            iWstb                                                  : in std_logic;
            oOverflow                                              : out std_logic;
            iOverflowClear                                         : in std_logic;
            oFifoPush                                              : out std_logic;
            oFifoDin                                               : out std_logic_vector(20 downto 0);
            iFifoFull                                              : in std_logic;
            iFifoOverFlow                                          : in std_logic;
            iEvents                                                : in IdefxEventVector_t
        );
    end component;
    component Calibration is 
        port (
            iClk                                                   : in std_logic;
            iRst_n                                                 : in std_logic;
            iWstb                                                  : in std_logic;
            iTq                                                    : in std_logic_vector(15 downto 0);
            iDmask                                                 : in std_logic_vector(31 downto 0);
            i15u2Tick                                              : in std_logic;
            iEvent                                                 : in std_logic_vector(20 downto 0);
            iIrq                                                   : in std_logic;
            i1msTick                                               : in std_logic;
            iSWClear                                               : in std_logic;
            iSWEn                                                  : in std_logic;
            oSWRdy                                                 : out std_logic;
            oSWIrq                                                 : out std_logic;
            oEnable                                                : out std_logic;
            oCounter                                               : out std_logic_vector(31 downto 0);
            oTruncate                                              : out std_logic_vector(20 downto 0)
        );
    end component;
    component Incrementer16 is 
        generic (
            Technology                                             : integer
        );
        port (
            DataA                                                  : in std_logic_vector(15 downto 0);
            Sum                                                    : out std_logic_vector(15 downto 0)
        );
    end component;
    component Incrementer24 is 
        generic (
            Technology                                             : integer
        );
        port (
            DataA                                                  : in std_logic_vector(23 downto 0);
            Sum                                                    : out std_logic_vector(23 downto 0)
        );
    end component;
    component SramWrap is 
        generic (
            Technology                                             : integer
        );
        port (
            iClk                                                   : in std_logic;
            iRst_n                                                 : in std_logic;
            iEnable                                                : in std_logic;
            oFsmAddr                                               : out std_logic_vector(8 downto 0);
            oFsmAdcVal                                             : out std_logic_vector(11 downto 0);
            oFsmAdcCorr                                            : out std_logic_vector(11 downto 0);
            oFsmEnergy                                             : out std_logic_vector(4 downto 0);
            oSramWr                                                : out std_logic;
            oSramRd                                                : out std_logic;
            iSramDout                                              : in std_logic_vector(31 downto 0);
            iSramReady                                             : in std_logic;
            oSramDin                                               : out std_logic_vector(31 downto 0);
            oSramAddr                                              : out std_logic_vector(18 downto 0);
            oBramTrigWr                                            : out std_logic;
            oBramTrigRd                                            : out std_logic;
            iBramTrigDout                                          : in std_logic_vector(23 downto 0);
            iBramTrigReady                                         : in std_logic;
            oBramTrigDin                                           : out std_logic_vector(23 downto 0);
            oBramTrigAddr                                          : out std_logic_vector(4 downto 0);
            oBram1Wr                                               : out std_logic;
            oBram1Rd                                               : out std_logic;
            iBram1Dout                                             : in std_logic_vector(15 downto 0);
            iBram1Ready                                            : in std_logic;
            oBram1Din                                              : out std_logic_vector(15 downto 0);
            oBram1Addr                                             : out std_logic_vector(7 downto 0);
            oBram4Wr                                               : out std_logic;
            oBram4Rd                                               : out std_logic;
            iBram4Dout                                             : in std_logic_vector(23 downto 0);
            iBram4Ready                                            : in std_logic;
            oBram4Din                                              : out std_logic_vector(23 downto 0);
            oBram4Addr                                             : out std_logic_vector(5 downto 0);
            oFifoPop                                               : out std_logic;
            iFifoPush                                              : in std_logic;
            iFifoDout                                              : in std_logic_vector(20 downto 0);
            iFifoEmpty                                             : in std_logic;
            iFifoFull                                              : in std_logic;
            iAccNumQl                                              : in std_logic_vector(5 downto 0);
            iActiveNominal                                         : in std_logic;
            iActiveQl                                              : in std_logic_vector(1 downto 0);
            iActiveTLut                                            : in std_logic;
            oCount                                                 : out std_logic;
            iQlVarEmask                                            : in std_logic_vector(31 downto 0);
            iQlVarDmask                                            : in std_logic_vector(31 downto 0);
            iQlVarPmask                                            : in std_logic_vector(11 downto 0);
            iSumEMask                                              : in std_logic_vector(31 downto 0);
            iSumDMask                                              : in std_logic_vector(31 downto 0);
            oCalib                                                 : out std_logic;
            oCalibEvent                                            : out std_logic_vector(20 downto 0)
        );
    end component;
    component EventCounter is 
        port (
            iClk                                                   : in std_logic;
            iRst_n                                                 : in std_logic;
            iEnable                                                : in std_logic;
            iClear                                                 : in std_logic;
            iCount                                                 : in std_logic;
            oEventCount                                            : out std_logic_vector(31 downto 0)
        );
    end component;
    component IntCounter is 
        port (
            iClk                                                   : in std_logic;
            iRst_n                                                 : in std_logic;
            iReset                                                 : in std_logic;
            iWstb                                                  : in std_logic;
            iSetEnable                                             : in std_logic;
            iClearEnable                                           : in std_logic;
            i100msTick                                             : in std_logic;
            iQlIntTime                                             : in std_logic_vector(15 downto 0);
            iQlClear                                               : in std_logic;
            iIntTimeMin                                            : in std_logic_vector(15 downto 0);
            iIntTimeMax                                            : in std_logic_vector(15 downto 0);
            iIntEventsMax                                          : in std_logic_vector(31 downto 0);
            iEventCount                                            : in std_logic_vector(31 downto 0);
            oEnable                                                : out std_logic;
            oQlReady                                               : out std_logic;
            oQlIrq                                                 : out std_logic;
            oReset                                                 : out std_logic;
            oEventClear                                            : out std_logic;
            oActiveNominal                                         : out std_logic;
            oActiveQl                                              : out std_logic_vector(1 downto 0);
            oAccNumQl                                              : out std_logic_vector(5 downto 0)
        );
    end component;
    component EdgeDetect is 
        port (
            async_sig                                              : in std_logic;
            clk                                                    : in std_logic;
            rise                                                   : out std_logic;
            fall                                                   : out std_logic;
            rst_n                                                  : in std_logic
        );
    end component;
    component PulseGen is 
        port (
            clk                                                    : in std_logic;
            rst_n                                                  : in std_logic;
            pulse_in                                               : in std_logic;
            pulse_out                                              : out std_logic
        );
    end component;
    component ReadoutFsm is 
        generic (
            Technology                                             : integer
        );
        port (
            iEvents                                                : in IdefxEventVector_t;
            iClk                                                   : in std_logic;
            iRst_n                                                 : in std_logic;
            iApb                                                   : in ReadoutFsmIn_t;
            oApb                                                   : out ReadoutFsmOut_t;
            iCache                                                 : in CacheDetOut_t;
            oCache                                                 : out CacheDetIn_t;
            oRotb                                                  : out RotbDetIn_t;
            i100msTick                                             : in std_logic;
            i1msTick                                               : in std_logic;
            i15u2Tick                                              : in std_logic
        );
    end component;
    component TestPulse is 
        port (
            iClk                                                   : in std_logic;
            iRst_n                                                 : in std_logic;
            iTestStb                                               : in std_logic;
            i15u2Tick                                              : in std_logic;
            oBusy                                                  : out std_logic;
            oTestPulse                                             : out std_logic;
            oDacGo                                                 : out std_logic;
            iDacIrq                                                : in std_logic
        );
    end component;
    component DacCtrl is 
        port (
            iClk                                                   : in std_logic;
            iRst_n                                                 : in std_logic;
            iDin                                                   : in std_logic_vector(11 downto 0);
            iMode                                                  : in std_logic_vector(1 downto 0);
            iGo                                                    : in std_logic;
            oIrq                                                   : out std_logic;
            i800nsTick                                             : in std_logic;
            oSclk                                                  : out std_logic;
            oDin                                                   : out std_logic;
            oSync_n                                                : out std_logic
        );
    end component;
    component QuarterCtrl is 
        generic (
            Technology                                             : integer
        );
        port (
            iRst_n                                                 : in std_logic;
            iQctrl                                                 : in QuarterCtrlIn_t;
            oQctrl                                                 : out QuarterCtrlOut_t;
            oQuarters                                              : out QuarterInVector_t;
            iQuarters                                              : in QuarterOutVector_t;
            iClk                                                   : in std_logic;
            i15u2Tick                                              : in std_logic;
            i800nsTick                                             : in std_logic
        );
    end component;
    component DetCtrl is 
        generic (
            Technology                                             : integer
        );
        port (
            iClkM                                                  : in std_logic;
            iRstM_n                                                : in std_logic;
            iCache                                                 : in CacheDetOut_t;
            oCache                                                 : out CacheDetIn_t;
            iApb                                                   : in ApbDetOut_t;
            oApb                                                   : out ApbDetIn_t;
            oRotb                                                  : out RotbDetIn_t;
            iPin                                                   : in DetPinIn_t;
            oPin                                                   : out DetPinOut_t;
            i100msTick                                             : in std_logic;
            iClkF                                                  : in std_logic;
            i1msTick                                               : in std_logic;
            i800nsTick                                             : in std_logic;
            i15u2Tick                                              : in std_logic;
            iRstF_n                                                : in std_logic
        );
    end component;
    component ApbWrap is 
        generic (
            pIndex                                                 : integer;
            pAddr                                                  : integer;
            pMask                                                  : integer;
            pIrq                                                   : integer;
            PROT_CHANNEL_NUMBER                                    : integer
        );
        port (
            iClk                                                   : in std_logic;
            iRst_n                                                 : in std_logic;
            oCache                                                 : out ApbCacheOut_t;
            iCache                                                 : in ApbCacheIn_t;
            oDet                                                   : out ApbDetOut_t;
            iDet                                                   : in ApbDetIn_t;
            oRotb                                                  : out ApbRotbOut_t;
            iRotb                                                  : in ApbRotbIn_t;
            iApb                                                   : in apb_slv_in_type;
            oApb                                                   : out apb_slv_out_type;
            iAs                                                    : in ApbAsIn_t;
            oAs                                                    : out ApbAsOut_t;
            iHk                                                    : in ApbHkIn_t;
            oHk                                                    : out ApbHkOut_t;
            iTimer                                                 : in ApbTimerIn_t;
            oTimer                                                 : out ApbTimerOut_t;
            iAttn                                                  : in ApbAttnIn_t;
            oAttn                                                  : out ApbAttnOut_t;
            iGenReg                                                : in ApbGenRegIn_t;
            oGenReg                                                : out ApbGenRegOut_t
        );
    end component;
    component PinWrap is 
        generic (
            StrobeInverted                                         : integer;
            Technology                                             : integer;
            AdcDoutInverted                                        : integer
        );
        port (
            iDet                                                   : in DetPinOut_t;
            oDet                                                   : out DetPinIn_t;
            iDetDout_n                                             : in std_logic_vector(1 to 16);
            iDetDout_p                                             : in std_logic_vector(1 to 16);
            oDetDin_n                                              : out std_logic_vector(1 to 16);
            oDetDin_p                                              : out std_logic_vector(1 to 16);
            oDetStrobe_n                                           : out std_logic_vector(1 to 16);
            oDetStrobe_p                                           : out std_logic_vector(1 to 16);
            iDetAdcDout                                            : in std_logic_vector(1 to 16);
            oDetAdcCs                                              : out std_logic_vector(1 to 16);
            oDetAdcSclk                                            : out std_logic_vector(1 to 16);
            oDetQDacDin                                            : out std_logic_vector(1 to 4);
            oDetQDacSclk                                           : out std_logic_vector(1 to 4);
            oDetQDacSync_n                                         : out std_logic_vector(1 to 4);
            oDetQOn                                                : out std_logic_vector(1 to 4);
            oDetQTestPulse                                         : out std_logic_vector(1 to 4);
            iDetQSeu                                               : in std_logic_vector(1 to 4);
            iEn                                                    : in std_logic;
            iClk                                                   : in std_logic
        );
    end component;
    component RotbSdWrap is 
        generic (
            USE_EDAC                                               : integer;
            USE_SCRUB                                              : integer
        );
        port (
            iAddr                                                  : in std_logic_vector(23 downto 0);
            iData                                                  : in std_logic_vector(31 downto 0);
            iEnable                                                : in std_logic;
            iRd                                                    : in std_logic;
            iRst_n                                                 : in std_logic;
            iSdq                                                   : in std_logic_vector(15 downto 0);
            iWr                                                    : in std_logic;
            oReady                                                 : out std_logic;
            oData                                                  : out std_logic_vector(31 downto 0);
            oDeDetected                                            : out std_logic;
            oInitialized                                           : out std_logic;
            oSa                                                    : out std_logic_vector(12 downto 0);
            oSba                                                   : out std_logic_vector(1 downto 0);
            oScas_n                                                : out std_logic;
            oScke                                                  : out std_logic;
            oSclk                                                  : out std_logic;
            oScs_n                                                 : out std_logic;
            oSdq                                                   : out std_logic_vector(15 downto 0);
            oSdqBdrive                                             : out std_logic;
            oSdqm                                                  : out std_logic_vector(1 downto 0);
            oSecCount                                              : out std_logic_vector(7 downto 0);
            oSras_n                                                : out std_logic;
            oSwe_n                                                 : out std_logic;
            iScrubRate                                             : in std_logic_vector(1 downto 0);
            iEdacOn                                                : in std_logic;
            iRefreshRate                                           : in std_logic_vector(7 downto 0);
            iEdacReset                                             : in std_logic;
            iClk                                                   : in std_logic;
            oAhb                                                   : out AhbRotbIn_t;
            iAhb                                                   : in AhbRotbOut_t;
            iCurrentBlock                                          : in std_logic_vector(16 downto 0);
            iCmdStrobe                                             : in std_logic;
            iTick15u2                                              : in std_logic;
            iTick800ns                                             : in std_logic;
            oIrq                                                   : out std_logic
        );
    end component;
    component RotbCtrl is 
        generic (
            MAX_BLOCKS                                             : integer;
            USE_EDAC                                               : integer;
            USE_SCRUB                                              : integer
        );
        port (
            iDet                                                   : in RotbDetIn_t;
            iClk                                                   : in std_logic;
            iRst_n                                                 : in std_logic;
            iApb                                                   : in ApbRotbOut_t;
            oApb                                                   : out ApbRotbIn_t;
            oROTBa                                                 : out std_logic_vector(12 downto 0);
            oROTBba                                                : out std_logic_vector(1 downto 0);
            oROTBdqm                                               : out std_logic_vector(1 downto 0);
            oROTBcke                                               : out std_logic;
            oROTBclk                                               : out std_logic;
            oROTBcs_n                                              : out std_logic;
            oROTBcas_n                                             : out std_logic;
            oROTBras_n                                             : out std_logic;
            oROTBwe_n                                              : out std_logic;
            oAs                                                    : out RotbAsOut_t;
            iAs                                                    : in RotbAsIn_t;
            iCache                                                 : in CacheRotbOut_t;
            oCache                                                 : out CacheRotbIn_t;
            oROTBdq                                                : out std_logic_vector(15 downto 0);
            oROTBdqBdrive                                          : out std_logic;
            iROTBdq                                                : in std_logic_vector(15 downto 0);
            iTimestamp                                             : in std_logic_vector(47 downto 0);
            iAhb                                                   : in AhbRotbOut_t;
            oAhb                                                   : out AhbRotbIn_t;
            iTick15u2                                              : in std_logic;
            iTick800ns                                             : in std_logic
        );
    end component;
    component HkAdcCtrl is 
        port (
            iADDR                                                  : in std_logic_vector(2 downto 0);
            iCLK                                                   : in std_logic;
            iGO                                                    : in std_logic;
            iRST_N                                                 : in std_logic;
            oCS_N                                                  : out std_logic;
            oDIN                                                   : out std_logic;
            oRDY                                                   : out std_logic;
            oSCLK                                                  : out std_logic;
            iDout                                                  : in std_logic;
            oDataVal                                               : out std_logic_vector(11 downto 0);
            iSclkTick                                              : in std_logic
        );
    end component;
    component hkmonitor is 
        generic (
            PROT_CHANNEL_NUMBER                                    : integer;
            UNLOCKING_TOKEN                                        : integer;
            TRACK_PRESCALER                                        : integer;
            DPU_1V5_C_MAX                                          : integer;
            DPU_2V5_C_MAX                                          : integer;
            DPU_3V3_C_MAX                                          : integer;
            DPU_SPW_C_MAX                                          : integer;
            DET_C_MAX                                              : integer;
            ATT_C_MAX                                              : integer;
            ATT_V_MAX                                              : integer;
            HV_01_V_MAX                                            : integer;
            HV_17_V_MAX                                            : integer
        );
        port (
            iAdcDout                                               : in std_logic;
            iClk                                                   : in std_logic;
            iRst_n                                                 : in std_logic;
            oAdcCs_n                                               : out std_logic_vector(1 to 2);
            oAdcDin                                                : out std_logic;
            oAdcSclk                                               : out std_logic;
            oMux                                                   : out std_logic_vector(1 downto 0);
            oAdcVal                                                : out std_logic_vector(11 downto 0);
            oIrq                                                   : out std_logic;
            oThresholds                                            : out HkThresholdVector_t;
            oProtStat                                              : out std_logic_vector(1 to 9);
            oProtEn                                                : out std_logic_vector(1 to 9);
            oAdcReady                                              : out std_logic;
            iProtEn                                                : in std_logic_vector(1 to 9);
            iIrqEn                                                 : in std_logic_vector(1 to 9);
            iAdcGo                                                 : in std_logic;
            iAdcAddress                                            : in std_logic_vector(5 downto 0);
            iToken                                                 : in std_logic_vector(7 downto 0);
            iTokenWrStb                                            : in std_logic;
            iThresholds                                            : in HkThresholdVector_t;
            iThreshWrStb                                           : in std_logic_vector(1 to 9);
            iProtClear                                             : in std_logic_vector(1 to 9);
            oBadSample                                             : out std_logic_vector(11 downto 0);
            i800nsTick                                             : in std_logic
        );
    end component;
    component ScanCtrl is 
        generic (
            Technology                                             : integer
        );
        port (
            oHkAdcAddress                                          : out std_logic_vector(5 downto 0);
            iHkAdcReady                                            : in std_logic;
            oHkAdcGo                                               : out std_logic;
            oAdcReady                                              : out std_logic;
            oAdcVal                                                : out std_logic_vector(11 downto 0);
            iHkAdcVal                                              : in std_logic_vector(11 downto 0);
            iAdcAddr                                               : in std_logic_vector(6 downto 0);
            oAsAdcGo                                               : out std_logic;
            oAsAdcAddress                                          : out std_logic_vector(3 downto 0);
            iAsAdcReady                                            : in std_logic_vector(1 downto 0);
            iAsAdcVal                                              : in std_logic_vector(11 downto 0);
            iClk                                                   : in std_logic;
            iRst_n                                                 : in std_logic
        );
    end component;
    component HkCtrl is 
        generic (
            PROT_CHANNEL_NUMBER                                    : integer;
            UNLOCKING_TOKEN                                        : integer;
            Technology                                             : integer;
            HV_LIMIT                                               : integer;
            DPU_1V5_C_MAX                                          : integer;
            DPU_2V5_C_MAX                                          : integer;
            DPU_3V3_C_MAX                                          : integer;
            DPU_SPW_C_MAX                                          : integer;
            DET_C_MAX                                              : integer;
            ATT_C_MAX                                              : integer;
            ATT_V_MAX                                              : integer;
            HV_01_V_MAX                                            : integer;
            HV_17_V_MAX                                            : integer;
            TRACK_PRESCALER                                        : integer
        );
        port (
            iRst_n                                                 : in std_logic;
            iClk                                                   : in std_logic;
            oApb                                                   : out ApbHkIn_t;
            iApb                                                   : in ApbHkOut_t;
            oAdcCs_n                                               : out std_logic_vector(1 to 2);
            oAdcDin                                                : out std_logic;
            iAdcDout                                               : in std_logic;
            oAdcSclk                                               : out std_logic;
            oPsuHvEnable                                           : out std_logic_vector(1 to 2);
            oPsuHvSet                                              : out std_logic_vector(1 to 2);
            oPsuLvEn                                               : out std_logic;
            oSpwEn                                                 : out std_logic_vector(1 downto 0);
            i800nsTick                                             : in std_logic;
            oAttnEn                                                : out std_logic;
            oMux                                                   : out std_logic_vector(1 downto 0);
            oDetEn                                                 : out std_logic;
            oAs                                                    : out AspHkIn_t;
            iAs                                                    : in AspHkOut_t
        );
    end component;
    component AsAdcCtrl is 
        port (
            iAddr                                                  : in std_logic_vector(2 downto 0);
            iClk                                                   : in std_logic;
            iGo                                                    : in std_logic;
            iRst_n                                                 : in std_logic;
            oCs_n                                                  : out std_logic;
            oDin                                                   : out std_logic;
            oRdy                                                   : out std_logic;
            oSclk                                                  : out std_logic;
            iDoutB                                                 : in std_logic;
            oDataValA                                              : out std_logic_vector(11 downto 0);
            iSclkTick                                              : in std_logic;
            iDoutA                                                 : in std_logic;
            oDataValB                                              : out std_logic_vector(11 downto 0)
        );
    end component;
    component AsCtrl is 
        generic (
            Technology                                             : integer;
            CsInverted                                             : integer
        );
        port (
            iRst_n                                                 : in std_logic;
            oApb                                                   : out ApbAsIn_t;
            iApb                                                   : in ApbAsOut_t;
            iClk                                                   : in std_logic;
            oASPaOn                                                : out std_logic;
            oASPaADCcs_n                                           : out std_logic;
            oASPaADCsclk                                           : out std_logic;
            oASPaADCdin                                            : out std_logic;
            iASPaADCdout                                           : in std_logic;
            oASPbOn                                                : out std_logic;
            oASPbADCcs_n                                           : out std_logic;
            oASPbADCsclk                                           : out std_logic;
            oASPbADCdin                                            : out std_logic;
            iASPbADCdout                                           : in std_logic;
            iRotb                                                  : in RotbAsOut_t;
            oRotb                                                  : out RotbAsIn_t;
            i1msTick                                               : in std_logic;
            iHk                                                    : in AspHkIn_t;
            oHk                                                    : out AspHkOut_t;
            iSclkTick                                              : in std_logic
        );
    end component;
    component LongTimer is 
        port (
            iRst_n                                                 : in std_logic;
            iClk                                                   : in std_logic;
            oApb                                                   : out ApbTimerIn_t;
            iApb                                                   : in ApbTimerOut_t;
            o100msTick                                             : out std_logic;
            o1msTick                                               : out std_logic;
            oTimestamp                                             : out std_logic_vector(47 downto 0);
            o800nsTick                                             : out std_logic;
            o15u2Tick                                              : out std_logic
        );
    end component;
    component attpwm is 
        port (
            iClk                                                   : in std_logic;
            iEna                                                   : in std_logic;
            ipwmDuty                                               : in std_logic_vector(8 downto 0);
            ipwmPeriod                                             : in std_logic_vector(7 downto 0);
            ipwmPrescale                                           : in std_logic_vector(3 downto 0);
            iRst_n                                                 : in std_logic;
            oPwmFallingEdge                                        : out std_logic;
            oPwmOutput                                             : out std_logic
        );
    end component;
    component AttnCtrl is 
        port (
            iRst_n                                                 : in std_logic;
            iClk                                                   : in std_logic;
            oApb                                                   : out ApbAttnIn_t;
            iApb                                                   : in ApbAttnOut_t;
            oAttnPwmA                                              : out std_logic;
            oAttnPwmB                                              : out std_logic;
            oAttnDirA                                              : out std_logic;
            oAttnDirB                                              : out std_logic;
            iAttnPosAb                                             : in std_logic;
            iAttnPosBc                                             : in std_logic;
            i10HzCE                                                : in std_logic;
            i1kHzCE                                                : in std_logic;
            iEn                                                    : in std_logic
        );
    end component;
    component SramCtrl is 
        generic (
            USE_EDAC                                               : integer
        );
        port (
            iClk                                                   : in std_logic;
            iRst_n                                                 : in std_logic;
            iEdacOn                                                : in std_logic;
            iWr                                                    : in std_logic;
            oSec                                                   : out std_logic;
            oReady                                                 : out std_logic;
            oData                                                  : out std_logic_vector(31 downto 0);
            iRd                                                    : in std_logic;
            iAddr                                                  : in std_logic_vector(18 downto 0);
            iData                                                  : in std_logic_vector(31 downto 0);
            oDed                                                   : out std_logic;
            oSramCe_n                                              : out std_logic_vector(3 downto 0);
            oSramWe_n                                              : out std_logic;
            oSramOe_n                                              : out std_logic;
            oSramBdrive                                            : out std_logic;
            oSramAddr                                              : out std_logic_vector(17 downto 0);
            oSramDout                                              : out std_logic_vector(31 downto 0);
            oSramCbout                                             : out std_logic_vector(6 downto 0);
            iSramDin                                               : in std_logic_vector(31 downto 0);
            iSramCbin                                              : in std_logic_vector(6 downto 0)
        );
    end component;
    component ScrubCtrl is 
        generic (
            ADDR_BIT                                               : integer
        );
        port (
            iClk                                                   : in std_logic;
            iRst_n                                                 : in std_logic;
            iTick15u2                                              : in std_logic;
            iTick800ns                                             : in std_logic;
            oRd                                                    : out std_logic;
            iScrubRate                                             : in std_logic_vector(1 downto 0);
            oAddr                                                  : out std_logic_vector(18 downto 0);
            iReady                                                 : in std_logic
        );
    end component;
    component CacheCtrl is 
        generic (
            Technology                                             : integer;
            USE_EDAC                                               : integer;
            USE_SCRUB                                              : integer
        );
        port (
            oDet                                                   : out CacheDetOut_t;
            iDet                                                   : in CacheDetIn_t;
            iClkm                                                  : in std_logic;
            iRstM_n                                                : in std_logic;
            iApb                                                   : in ApbCacheOut_t;
            oApb                                                   : out ApbCacheIn_t;
            oCACHEa                                                : out std_logic_vector(17 downto 0);
            iCACHEdq                                               : in std_logic_vector(31 downto 0);
            iCacheCb                                               : in std_logic_vector(6 downto 0);
            oCACHEwe_n                                             : out std_logic_vector(3 downto 0);
            oCACHEoe_n                                             : out std_logic_vector(3 downto 0);
            oCACHEce_n                                             : out std_logic_vector(3 downto 0);
            iClkf                                                  : in std_logic;
            oRotb                                                  : out CacheRotbOut_t;
            iRotb                                                  : in CacheRotbIn_t;
            oCACHEdq                                               : out std_logic_vector(31 downto 0);
            oCACHEdqBdrive                                         : out std_logic;
            oCacheCb                                               : out std_logic_vector(6 downto 0);
            oCACHEcbBdrive                                         : out std_logic;
            oAhb                                                   : out AhbCacheIn_t;
            iAhb                                                   : in AhbCacheOut_t;
            iTick800ns                                             : in std_logic;
            iTick15u2                                              : in std_logic;
            iRstF_n                                                : in std_logic
        );
    end component;
    component GenReg is 
        generic (
            SYSTEM_RELEASE                                         : integer;
            SYSTEM_BUILD                                           : integer;
            Technology                                             : integer;
            WDOG_RELOAD                                            : integer;
            WDOG_DISABLED                                          : integer;
            WDOG_PRESCALER                                         : integer
        );
        port (
            iRst_n                                                 : in std_logic;
            iClk                                                   : in std_logic;
            oApb                                                   : out ApbGenRegIn_t;
            iApb                                                   : in ApbGenRegOut_t;
            iOtherIdpuIsOn                                         : in std_logic;
            iThisIsMain                                            : in std_logic;
            oWatchDog                                              : out std_logic;
            oUseEeprom                                             : out std_logic;
            oTxTick                                                : out std_logic
        );
    end component;
    component AhbWrap is 
        generic (
            hIndex                                                 : integer;
            hAddr                                                  : integer;
            hMask                                                  : integer
        );
        port (
            iClk                                                   : in std_logic;
            iRst_n                                                 : in std_logic;
            oCache                                                 : out AhbCacheOut_t;
            iCache                                                 : in AhbCacheIn_t;
            oRotb                                                  : out AhbRotbOut_t;
            iRotb                                                  : in AhbRotbIn_t;
            iAhb                                                   : in ahb_slv_in_type;
            oAhb                                                   : out ahb_slv_out_type
        );
    end component;
    component StixCtrl is 
        generic (
            pAddr                                                  : integer;
            hIndex                                                 : integer;
            pIndex                                                 : integer;
            hAddr                                                  : integer;
            hMask                                                  : integer;
            pMask                                                  : integer;
            pIrq                                                   : integer;
            SYSTEM_RELEASE                                         : integer;
            SYSTEM_BUILD                                           : integer;
            Technology                                             : integer;
            PROT_CHANNEL_NUMBER                                    : integer;
            UNLOCKING_TOKEN                                        : integer;
            ROTB_MAX_BLOCKS                                        : integer;
            WDOG_RELOAD                                            : integer;
            WDOG_DISABLED                                          : integer;
            WDOG_PRESCALER                                         : integer;
            ROTB_EDAC_USE                                          : integer;
            ROTB_SCRUB_USE                                         : integer;
            CACHE_EDAC_USE                                         : integer;
            CACHE_SCRUB_USE                                        : integer;
            HV_LIMIT                                               : integer;
            TRACK_PRESCALER                                        : integer;
            DPU_1V5_C_MAX                                          : integer;
            DPU_2V5_C_MAX                                          : integer;
            DPU_3V3_C_MAX                                          : integer;
            DPU_SPW_C_MAX                                          : integer;
            DET_C_MAX                                              : integer;
            ATT_C_MAX                                              : integer;
            ATT_V_MAX                                              : integer;
            HV_01_V_MAX                                            : integer;
            HV_17_V_MAX                                            : integer
        );
        port (
            iRstM_n                                                : in std_logic;
            iClkm                                                  : in std_logic;
            iClkf                                                  : in std_logic;
            iApb                                                   : in apb_slv_in_type;
            oApb                                                   : out apb_slv_out_type;
            oROTBclk                                               : out std_logic;
            oROTBcke                                               : out std_logic;
            oROTBwe_n                                              : out std_logic;
            oROTBcas_n                                             : out std_logic;
            oROTBcs_n                                              : out std_logic;
            oROTBras_n                                             : out std_logic;
            iROTBdq                                                : in std_logic_vector(15 downto 0);
            oROTBa                                                 : out std_logic_vector(12 downto 0);
            oROTBba                                                : out std_logic_vector(1 downto 0);
            oROTBdqm                                               : out std_logic_vector(1 downto 0);
            oASPaOn                                                : out std_logic;
            oASPaADCcs_n                                           : out std_logic;
            oASPaADCsclk                                           : out std_logic;
            oASPaADCdin                                            : out std_logic;
            iASPaADCdout                                           : in std_logic;
            oASPbOn                                                : out std_logic;
            oASPbADCcs_n                                           : out std_logic;
            oASPbADCsclk                                           : out std_logic;
            oASPbADCdin                                            : out std_logic;
            iASPbADCdout                                           : in std_logic;
            oCACHEa                                                : out std_logic_vector(17 downto 0);
            iDetDout_n                                             : in std_logic_vector(1 to 16);
            iDetDout_p                                             : in std_logic_vector(1 to 16);
            oDetDin_n                                              : out std_logic_vector(1 to 16);
            oDetDin_p                                              : out std_logic_vector(1 to 16);
            oDetStrobe_n                                           : out std_logic_vector(1 to 16);
            oDetStrobe_p                                           : out std_logic_vector(1 to 16);
            iDetAdcDout                                            : in std_logic_vector(1 to 16);
            oDetAdcCs                                              : out std_logic_vector(1 to 16);
            oDetAdcSclk                                            : out std_logic_vector(1 to 16);
            oDetQDacDin                                            : out std_logic_vector(1 to 4);
            oDetQDacSclk                                           : out std_logic_vector(1 to 4);
            oDetQDacSync_n                                         : out std_logic_vector(1 to 4);
            oDetQOn                                                : out std_logic_vector(1 to 4);
            oDetQTestPulse                                         : out std_logic_vector(1 to 4);
            iDetQSeu                                               : in std_logic_vector(1 to 4);
            oAttnPwmA                                              : out std_logic;
            oAttnPwmB                                              : out std_logic;
            oAttnDirA                                              : out std_logic;
            oAttnDirB                                              : out std_logic;
            iAttnPosAb                                             : in std_logic;
            iAttnPosBc                                             : in std_logic;
            oPsuHvSet                                              : out std_logic_vector(1 to 2);
            oPsuLvEn                                               : out std_logic;
            oSpwEn                                                 : out std_logic_vector(1 downto 0);
            iOtherIdpuIsOn                                         : in std_logic;
            iThisIsMain                                            : in std_logic;
            oAhb                                                   : out ahb_slv_out_type;
            iAhb                                                   : in ahb_slv_in_type;
            oPsuHvEn                                               : out std_logic_vector(1 to 2);
            oAdcCs_n                                               : out std_logic_vector(1 to 2);
            oAdcDin                                                : out std_logic;
            iAdcDout                                               : in std_logic;
            oAdcSclk                                               : out std_logic;
            oCACHEwe_n                                             : out std_logic_vector(3 downto 0);
            oCACHEoe_n                                             : out std_logic_vector(3 downto 0);
            oCACHEce_n                                             : out std_logic_vector(3 downto 0);
            oROTBdq                                                : out std_logic_vector(15 downto 0);
            oROTBdqBdrive                                          : out std_logic;
            oCACHEdq                                               : out std_logic_vector(31 downto 0);
            oCACHEdqBdrive                                         : out std_logic;
            iCACHEdq                                               : in std_logic_vector(31 downto 0);
            iCacheCb                                               : in std_logic_vector(6 downto 0);
            oCacheCb                                               : out std_logic_vector(6 downto 0);
            oCACHEcbBdrive                                         : out std_logic;
            oUseEeprom                                             : out std_logic;
            oHkMux                                                 : out std_logic_vector(1 downto 0);
            oWatchDog                                              : out std_logic;
            oTick15u2                                              : out std_logic;
            oTick800ns                                             : out std_logic;
            oTick1ms                                               : out std_logic;
            iRstF_n                                                : in std_logic;
            oTxTick                                                : out std_logic;
            oTick100ms                                             : out std_logic;
            iClkFF                                                 : in std_logic
        );
    end component;
    component StixSpw is 
        generic (
            SysFreq                                                : integer;
            FabTech                                                : integer;
            MemTech                                                : integer;
            DestKey                                                : integer;
            NodeAddr                                               : integer;
            hIndex                                                 : integer;
            pIndex                                                 : integer;
            pIrq                                                   : integer;
            pMask                                                  : integer;
            pAddr                                                  : integer
        );
        port (
            iDat0                                                  : in std_logic;
            iStb0                                                  : in std_logic;
            oDat0                                                  : out std_logic;
            oStb0                                                  : out std_logic;
            oAhb                                                   : out ahb_mst_out_type;
            iAhb                                                   : in ahb_mst_in_type;
            iApb                                                   : in apb_slv_in_type;
            oApb                                                   : out apb_slv_out_type;
            iRst_n                                                 : in std_logic;
            iClk                                                   : in std_logic;
            iDat1                                                  : in std_logic;
            iStb1                                                  : in std_logic;
            oDat1                                                  : out std_logic;
            oStb1                                                  : out std_logic;
            iSpwEn                                                 : in std_logic_vector(1 downto 0)
        );
    end component;
    component StixRstGen is 
        generic (
            Technology                                             : integer
        );
        port (
            iClk                                                   : in std_logic;
            iClkM                                                  : in std_logic;
            iClkF                                                  : in std_logic;
            iExtRst_n                                              : in std_logic;
            iWdg                                                   : in std_logic;
            oRstM_n                                                : out std_logic;
            oRstF_n                                                : out std_logic;
            oRstFF_n                                               : out std_logic
        );
    end component;
    component StixIdpu is 
        generic (
            SYSTEM_RELEASE                                         : integer;
            SYSTEM_BUILD                                           : integer;
            Technology                                             : integer;
            UseEepromTypeBit                                       : integer
        );
        port (
            oConsoleTx                                             : out std_logic;
            iConsoleRx                                             : in std_logic;
            iJtagTck                                               : in std_logic;
            iJtagTms                                               : in std_logic;
            iJtagTdi                                               : in std_logic;
            oJtagTdo                                               : out std_logic;
            iSpw0Dat                                               : in std_logic;
            iSpw0Stb                                               : in std_logic;
            oSpw0Dat                                               : out std_logic;
            oSpw0Stb                                               : out std_logic;
            oRomCe_n                                               : out std_logic_vector(7 downto 0);
            iFbsy_n                                                : in std_logic_vector(1 to 2);
            oFale                                                  : out std_logic_vector(1 to 2);
            oFCe_n                                                 : out std_logic_vector(15 downto 0);
            oFcle                                                  : out std_logic_vector(1 to 2);
            oFre_n                                                 : out std_logic_vector(1 to 2);
            oFwe_n                                                 : out std_logic_vector(1 to 2);
            oFwp_n                                                 : out std_logic_vector(1 to 2);
            oDetDin_n                                              : out std_logic_vector(1 to 16);
            oDetDin_p                                              : out std_logic_vector(1 to 16);
            oDetStrobe_n                                           : out std_logic_vector(1 to 16);
            oDetStrobe_p                                           : out std_logic_vector(1 to 16);
            iDetDout_n                                             : in std_logic_vector(1 to 16);
            iDetDout_p                                             : in std_logic_vector(1 to 16);
            oDetAdcCs                                              : out std_logic_vector(1 to 16);
            oDetAdcSclk                                            : out std_logic_vector(1 to 16);
            iDetAdcDout                                            : in std_logic_vector(1 to 16);
            oDetQDacSync_n                                         : out std_logic_vector(1 to 4);
            oDetQDacSclk                                           : out std_logic_vector(1 to 4);
            oDetQDacDin                                            : out std_logic_vector(1 to 4);
            oDetQOn                                                : out std_logic_vector(1 to 4);
            oDetQTestPulse                                         : out std_logic_vector(1 to 4);
            iDetQSeu                                               : in std_logic_vector(1 to 4);
            oASPaOn                                                : out std_logic;
            oASPaADCcs_n                                           : out std_logic;
            oASPaADCsclk                                           : out std_logic;
            oASPaADCdin                                            : out std_logic;
            iASPaADCdout                                           : in std_logic;
            oASPbOn                                                : out std_logic;
            oASPbADCcs_n                                           : out std_logic;
            oASPbADCsclk                                           : out std_logic;
            oASPbADCdin                                            : out std_logic;
            iASPbADCdout                                           : in std_logic;
            oCACHEa                                                : out std_logic_vector(17 downto 0);
            oPsuHvEn                                               : out std_logic_vector(1 to 2);
            oPsuHvSet                                              : out std_logic_vector(1 to 2);
            oPsuLvEn                                               : out std_logic;
            oAttnPwmA                                              : out std_logic;
            oAttnPwmB                                              : out std_logic;
            oAttnDirA                                              : out std_logic;
            oAttnDirB                                              : out std_logic;
            iAttnPosAb                                             : in std_logic;
            iAttnPosBc                                             : in std_logic;
            iOtherIdpuIsOn                                         : in std_logic;
            iThisIsMain                                            : in std_logic;
            iSpw1Dat                                               : in std_logic;
            iSpw1Stb                                               : in std_logic;
            oSpw1Dat                                               : out std_logic;
            oSpw1Stb                                               : out std_logic;
            iExtRst_n                                              : in std_logic;
            iClk                                                   : in std_logic;
            oR2clk                                                 : out std_logic;
            oR2cke                                                 : out std_logic;
            oR2ba                                                  : out std_logic_vector(1 downto 0);
            oR1clk                                                 : out std_logic;
            oR1cke                                                 : out std_logic;
            oR1ba                                                  : out std_logic_vector(1 downto 0);
            oR2a                                                   : out std_logic_vector(12 downto 0);
            oR1a                                                   : out std_logic_vector(12 downto 0);
            oR1dqm                                                 : out std_logic_vector(1 downto 0);
            oR2dqm                                                 : out std_logic_vector(1 downto 0);
            oR2cs_n                                                : out std_logic;
            oR1cs_n                                                : out std_logic;
            oR2we_n                                                : out std_logic;
            oR1we_n                                                : out std_logic;
            oR2cas_n                                               : out std_logic;
            oR1cas_n                                               : out std_logic;
            oR2ras_n                                               : out std_logic;
            oR1ras_n                                               : out std_logic;
            oAdcCs_n                                               : out std_logic_vector(1 to 2);
            oAdcDin                                                : out std_logic;
            iAdcDout                                               : in std_logic;
            oAdcSclk                                               : out std_logic;
            oCACHEwe_n                                             : out std_logic_vector(3 downto 0);
            oCACHEoe_n                                             : out std_logic_vector(3 downto 0);
            oCACHEce_n                                             : out std_logic_vector(3 downto 0);
            iRomBsy_n                                              : in std_logic;
            oRomRst_n                                              : out std_logic;
            oRomOe_n                                               : out std_logic;
            oRomWe_n                                               : out std_logic;
            oRomA                                                  : out std_logic_vector(16 downto 0);
            iCACHEdq                                               : in std_logic_vector(31 downto 0);
            oCACHEdq                                               : out std_logic_vector(31 downto 0);
            oCACHEdqBdrive                                         : out std_logic;
            oCACHEcbBdrive                                         : out std_logic;
            oRomIoBdrive                                           : out std_logic;
            iRomIo                                                 : in std_logic_vector(7 downto 0);
            oRomIo                                                 : out std_logic_vector(7 downto 0);
            iFio                                                   : in std_logic_vector(15 downto 0);
            oFio                                                   : out std_logic_vector(15 downto 0);
            oFioBdrive                                             : out std_logic;
            oUseEeprom                                             : out std_logic;
            oR1dq                                                  : out std_logic_vector(15 downto 0);
            oR1dqBdrive                                            : out std_logic;
            oR2dqBdrive                                            : out std_logic;
            oR2dq                                                  : out std_logic_vector(15 downto 0);
            iR1dq                                                  : in std_logic_vector(15 downto 0);
            iR2dq                                                  : in std_logic_vector(15 downto 0);
            oHkMux                                                 : out std_logic_vector(1 downto 0);
            iCacheCb                                               : in std_logic_vector(6 downto 0);
            oCacheCb                                               : out std_logic_vector(6 downto 0);
            oSpwEn                                                 : out std_logic_vector(1 to 2)
        );
    end component;
end package Stix_pkg;
